//Generate the verilog at 2025-10-17T18:45:31 by iSTA.
module top (
clk,
reset,
alu_result_out,
load_data_out,
pc_out
);

input clk ;
input reset ;
output [31:0] alu_result_out ;
output [31:0] load_data_out ;
output [31:0] pc_out ;

wire _00000_ ;
wire _00001_ ;
wire _00002_ ;
wire _00003_ ;
wire _00004_ ;
wire _00005_ ;
wire _00006_ ;
wire _00007_ ;
wire _00008_ ;
wire _00009_ ;
wire _00010_ ;
wire _00011_ ;
wire _00012_ ;
wire _00013_ ;
wire _00014_ ;
wire _00015_ ;
wire _00016_ ;
wire _00017_ ;
wire _00018_ ;
wire _00019_ ;
wire _00020_ ;
wire _00021_ ;
wire _00022_ ;
wire _00023_ ;
wire _00024_ ;
wire _00025_ ;
wire _00026_ ;
wire _00027_ ;
wire _00028_ ;
wire _00029_ ;
wire _00030_ ;
wire _00031_ ;
wire _00032_ ;
wire _00033_ ;
wire _00034_ ;
wire _00035_ ;
wire _00036_ ;
wire _00037_ ;
wire _00038_ ;
wire _00039_ ;
wire _00040_ ;
wire _00041_ ;
wire _00042_ ;
wire _00043_ ;
wire _00044_ ;
wire _00045_ ;
wire _00046_ ;
wire _00047_ ;
wire _00048_ ;
wire _00049_ ;
wire _00050_ ;
wire _00051_ ;
wire _00052_ ;
wire _00053_ ;
wire _00054_ ;
wire _00055_ ;
wire _00056_ ;
wire _00057_ ;
wire _00058_ ;
wire _00059_ ;
wire _00060_ ;
wire _00061_ ;
wire _00062_ ;
wire _00063_ ;
wire _00064_ ;
wire _00065_ ;
wire _00066_ ;
wire _00067_ ;
wire _00068_ ;
wire _00069_ ;
wire _00070_ ;
wire _00071_ ;
wire _00072_ ;
wire _00073_ ;
wire _00074_ ;
wire _00075_ ;
wire _00076_ ;
wire _00077_ ;
wire _00078_ ;
wire _00079_ ;
wire _00080_ ;
wire _00081_ ;
wire _00082_ ;
wire _00083_ ;
wire _00084_ ;
wire _00085_ ;
wire _00086_ ;
wire _00087_ ;
wire _00088_ ;
wire _00089_ ;
wire _00090_ ;
wire _00091_ ;
wire _00092_ ;
wire _00093_ ;
wire _00094_ ;
wire _00095_ ;
wire _00096_ ;
wire _00097_ ;
wire _00098_ ;
wire _00099_ ;
wire _00100_ ;
wire _00101_ ;
wire _00102_ ;
wire _00103_ ;
wire _00104_ ;
wire _00105_ ;
wire _00106_ ;
wire _00107_ ;
wire _00108_ ;
wire _00109_ ;
wire _00110_ ;
wire _00111_ ;
wire _00112_ ;
wire _00113_ ;
wire _00114_ ;
wire _00115_ ;
wire _00116_ ;
wire _00117_ ;
wire _00118_ ;
wire _00119_ ;
wire _00120_ ;
wire _00121_ ;
wire _00122_ ;
wire _00123_ ;
wire _00124_ ;
wire _00125_ ;
wire _00126_ ;
wire _00127_ ;
wire _00128_ ;
wire _00129_ ;
wire _00130_ ;
wire _00131_ ;
wire _00132_ ;
wire _00133_ ;
wire _00134_ ;
wire _00135_ ;
wire _00136_ ;
wire _00137_ ;
wire _00138_ ;
wire _00139_ ;
wire _00140_ ;
wire _00141_ ;
wire _00142_ ;
wire _00143_ ;
wire _00144_ ;
wire _00145_ ;
wire _00146_ ;
wire _00147_ ;
wire _00148_ ;
wire _00149_ ;
wire _00150_ ;
wire _00151_ ;
wire _00152_ ;
wire _00153_ ;
wire _00154_ ;
wire _00155_ ;
wire _00156_ ;
wire _00157_ ;
wire _00158_ ;
wire _00159_ ;
wire _00160_ ;
wire _00161_ ;
wire _00162_ ;
wire _00163_ ;
wire _00164_ ;
wire _00165_ ;
wire _00166_ ;
wire _00167_ ;
wire _00168_ ;
wire _00169_ ;
wire _00170_ ;
wire _00171_ ;
wire _00172_ ;
wire _00173_ ;
wire _00174_ ;
wire _00175_ ;
wire _00176_ ;
wire _00177_ ;
wire _00178_ ;
wire _00179_ ;
wire _00180_ ;
wire _00181_ ;
wire _00182_ ;
wire _00183_ ;
wire _00184_ ;
wire _00185_ ;
wire _00186_ ;
wire _00187_ ;
wire _00188_ ;
wire _00189_ ;
wire _00190_ ;
wire _00191_ ;
wire _00192_ ;
wire _00193_ ;
wire _00194_ ;
wire _00195_ ;
wire _00196_ ;
wire _00197_ ;
wire _00198_ ;
wire _00199_ ;
wire _00200_ ;
wire _00201_ ;
wire _00202_ ;
wire _00203_ ;
wire _00204_ ;
wire _00205_ ;
wire _00206_ ;
wire _00207_ ;
wire _00208_ ;
wire _00209_ ;
wire _00210_ ;
wire _00211_ ;
wire _00212_ ;
wire _00213_ ;
wire _00214_ ;
wire _00215_ ;
wire _00216_ ;
wire _00217_ ;
wire _00218_ ;
wire _00219_ ;
wire _00220_ ;
wire _00221_ ;
wire _00222_ ;
wire _00223_ ;
wire _00224_ ;
wire _00225_ ;
wire _00226_ ;
wire _00227_ ;
wire _00228_ ;
wire _00229_ ;
wire _00230_ ;
wire _00231_ ;
wire _00232_ ;
wire _00233_ ;
wire _00234_ ;
wire _00235_ ;
wire _00236_ ;
wire _00237_ ;
wire _00238_ ;
wire _00239_ ;
wire _00240_ ;
wire _00241_ ;
wire _00242_ ;
wire _00243_ ;
wire _00244_ ;
wire _00245_ ;
wire _00246_ ;
wire _00247_ ;
wire _00248_ ;
wire _00249_ ;
wire _00250_ ;
wire _00251_ ;
wire _00252_ ;
wire _00253_ ;
wire _00254_ ;
wire _00255_ ;
wire _00256_ ;
wire _00257_ ;
wire _00258_ ;
wire _00259_ ;
wire _00260_ ;
wire _00261_ ;
wire _00262_ ;
wire _00263_ ;
wire _00264_ ;
wire _00265_ ;
wire _00266_ ;
wire _00267_ ;
wire _00268_ ;
wire _00269_ ;
wire _00270_ ;
wire _00271_ ;
wire _00272_ ;
wire _00273_ ;
wire _00274_ ;
wire _00275_ ;
wire _00276_ ;
wire _00277_ ;
wire _00278_ ;
wire _00279_ ;
wire _00280_ ;
wire _00281_ ;
wire _00282_ ;
wire _00283_ ;
wire _00284_ ;
wire _00285_ ;
wire _00286_ ;
wire _00287_ ;
wire _00288_ ;
wire _00289_ ;
wire _00290_ ;
wire _00291_ ;
wire _00292_ ;
wire _00293_ ;
wire _00294_ ;
wire _00295_ ;
wire _00296_ ;
wire _00297_ ;
wire _00298_ ;
wire _00299_ ;
wire _00300_ ;
wire _00301_ ;
wire _00302_ ;
wire _00303_ ;
wire _00304_ ;
wire _00305_ ;
wire _00306_ ;
wire _00307_ ;
wire _00308_ ;
wire _00309_ ;
wire _00310_ ;
wire _00311_ ;
wire _00312_ ;
wire _00313_ ;
wire _00314_ ;
wire _00315_ ;
wire _00316_ ;
wire _00317_ ;
wire _00318_ ;
wire _00319_ ;
wire _00320_ ;
wire _00321_ ;
wire _00322_ ;
wire _00323_ ;
wire _00324_ ;
wire _00325_ ;
wire _00326_ ;
wire _00327_ ;
wire _00328_ ;
wire _00329_ ;
wire _00330_ ;
wire _00331_ ;
wire _00332_ ;
wire _00333_ ;
wire _00334_ ;
wire _00335_ ;
wire _00336_ ;
wire _00337_ ;
wire _00338_ ;
wire _00339_ ;
wire _00340_ ;
wire _00341_ ;
wire _00342_ ;
wire _00343_ ;
wire _00344_ ;
wire _00345_ ;
wire _00346_ ;
wire _00347_ ;
wire _00348_ ;
wire _00349_ ;
wire _00350_ ;
wire _00351_ ;
wire _00352_ ;
wire _00353_ ;
wire _00354_ ;
wire _00355_ ;
wire _00356_ ;
wire _00357_ ;
wire _00358_ ;
wire _00359_ ;
wire _00360_ ;
wire _00361_ ;
wire _00362_ ;
wire _00363_ ;
wire _00364_ ;
wire _00365_ ;
wire _00366_ ;
wire _00367_ ;
wire _00368_ ;
wire _00369_ ;
wire _00370_ ;
wire _00371_ ;
wire _00372_ ;
wire _00373_ ;
wire _00374_ ;
wire _00375_ ;
wire _00376_ ;
wire _00377_ ;
wire _00378_ ;
wire _00379_ ;
wire _00380_ ;
wire _00381_ ;
wire _00382_ ;
wire _00383_ ;
wire _00384_ ;
wire _00385_ ;
wire _00386_ ;
wire _00387_ ;
wire _00388_ ;
wire _00389_ ;
wire _00390_ ;
wire _00391_ ;
wire _00392_ ;
wire _00393_ ;
wire _00394_ ;
wire _00395_ ;
wire _00396_ ;
wire _00397_ ;
wire _00398_ ;
wire _00399_ ;
wire _00400_ ;
wire _00401_ ;
wire _00402_ ;
wire _00403_ ;
wire _00404_ ;
wire _00405_ ;
wire _00406_ ;
wire _00407_ ;
wire _00408_ ;
wire _00409_ ;
wire _00410_ ;
wire _00411_ ;
wire _00412_ ;
wire _00413_ ;
wire _00414_ ;
wire _00415_ ;
wire _00416_ ;
wire _00417_ ;
wire _00418_ ;
wire _00419_ ;
wire _00420_ ;
wire _00421_ ;
wire _00422_ ;
wire _00423_ ;
wire _00424_ ;
wire _00425_ ;
wire _00426_ ;
wire _00427_ ;
wire _00428_ ;
wire _00429_ ;
wire _00430_ ;
wire _00431_ ;
wire _00432_ ;
wire _00433_ ;
wire _00434_ ;
wire _00435_ ;
wire _00436_ ;
wire _00437_ ;
wire _00438_ ;
wire _00439_ ;
wire _00440_ ;
wire _00441_ ;
wire _00442_ ;
wire _00443_ ;
wire _00444_ ;
wire _00445_ ;
wire _00446_ ;
wire _00447_ ;
wire _00448_ ;
wire _00449_ ;
wire _00450_ ;
wire _00451_ ;
wire _00452_ ;
wire _00453_ ;
wire _00454_ ;
wire _00455_ ;
wire _00456_ ;
wire _00457_ ;
wire _00458_ ;
wire _00459_ ;
wire _00460_ ;
wire _00461_ ;
wire _00462_ ;
wire _00463_ ;
wire _00464_ ;
wire _00465_ ;
wire _00466_ ;
wire _00467_ ;
wire _00468_ ;
wire _00469_ ;
wire _00470_ ;
wire _00471_ ;
wire _00472_ ;
wire _00473_ ;
wire _00474_ ;
wire _00475_ ;
wire _00476_ ;
wire _00477_ ;
wire _00478_ ;
wire _00479_ ;
wire _00480_ ;
wire _00481_ ;
wire _00482_ ;
wire _00483_ ;
wire _00484_ ;
wire _00485_ ;
wire _00486_ ;
wire _00487_ ;
wire _00488_ ;
wire _00489_ ;
wire _00490_ ;
wire _00491_ ;
wire _00492_ ;
wire _00493_ ;
wire _00494_ ;
wire _00495_ ;
wire _00496_ ;
wire _00497_ ;
wire _00498_ ;
wire _00499_ ;
wire _00500_ ;
wire _00501_ ;
wire _00502_ ;
wire _00503_ ;
wire _00504_ ;
wire _00505_ ;
wire _00506_ ;
wire _00507_ ;
wire _00508_ ;
wire _00509_ ;
wire _00510_ ;
wire _00511_ ;
wire _00512_ ;
wire _00513_ ;
wire _00514_ ;
wire _00515_ ;
wire _00516_ ;
wire _00517_ ;
wire _00518_ ;
wire _00519_ ;
wire _00520_ ;
wire _00521_ ;
wire _00522_ ;
wire _00523_ ;
wire _00524_ ;
wire _00525_ ;
wire _00526_ ;
wire _00527_ ;
wire _00528_ ;
wire _00529_ ;
wire _00530_ ;
wire _00531_ ;
wire _00532_ ;
wire _00533_ ;
wire _00534_ ;
wire _00535_ ;
wire _00536_ ;
wire _00537_ ;
wire _00538_ ;
wire _00539_ ;
wire _00540_ ;
wire _00541_ ;
wire _00542_ ;
wire _00543_ ;
wire _00544_ ;
wire _00545_ ;
wire _00546_ ;
wire _00547_ ;
wire _00548_ ;
wire _00549_ ;
wire _00550_ ;
wire _00551_ ;
wire _00552_ ;
wire _00553_ ;
wire _00554_ ;
wire _00555_ ;
wire _00556_ ;
wire _00557_ ;
wire _00558_ ;
wire _00559_ ;
wire _00560_ ;
wire _00561_ ;
wire _00562_ ;
wire _00563_ ;
wire _00564_ ;
wire _00565_ ;
wire _00566_ ;
wire _00567_ ;
wire _00568_ ;
wire _00569_ ;
wire _00570_ ;
wire _00571_ ;
wire _00572_ ;
wire _00573_ ;
wire _00574_ ;
wire _00575_ ;
wire _00576_ ;
wire _00577_ ;
wire _00578_ ;
wire _00579_ ;
wire _00580_ ;
wire _00581_ ;
wire _00582_ ;
wire _00583_ ;
wire _00584_ ;
wire _00585_ ;
wire _00586_ ;
wire _00587_ ;
wire _00588_ ;
wire _00589_ ;
wire _00590_ ;
wire _00591_ ;
wire _00592_ ;
wire _00593_ ;
wire _00594_ ;
wire _00595_ ;
wire _00596_ ;
wire _00597_ ;
wire _00598_ ;
wire _00599_ ;
wire _00600_ ;
wire _00601_ ;
wire _00602_ ;
wire _00603_ ;
wire _00604_ ;
wire _00605_ ;
wire _00606_ ;
wire _00607_ ;
wire _00608_ ;
wire _00609_ ;
wire _00610_ ;
wire _00611_ ;
wire _00612_ ;
wire _00613_ ;
wire _00614_ ;
wire _00615_ ;
wire _00616_ ;
wire _00617_ ;
wire _00618_ ;
wire _00619_ ;
wire _00620_ ;
wire _00621_ ;
wire _00622_ ;
wire _00623_ ;
wire _00624_ ;
wire _00625_ ;
wire _00626_ ;
wire _00627_ ;
wire _00628_ ;
wire _00629_ ;
wire _00630_ ;
wire _00631_ ;
wire _00632_ ;
wire _00633_ ;
wire _00634_ ;
wire _00635_ ;
wire _00636_ ;
wire _00637_ ;
wire _00638_ ;
wire _00639_ ;
wire _00640_ ;
wire _00641_ ;
wire _00642_ ;
wire _00643_ ;
wire _00644_ ;
wire _00645_ ;
wire _00646_ ;
wire _00647_ ;
wire _00648_ ;
wire _00649_ ;
wire _00650_ ;
wire _00651_ ;
wire _00652_ ;
wire _00653_ ;
wire _00654_ ;
wire _00655_ ;
wire _00656_ ;
wire _00657_ ;
wire _00658_ ;
wire _00659_ ;
wire _00660_ ;
wire _00661_ ;
wire _00662_ ;
wire _00663_ ;
wire _00664_ ;
wire _00665_ ;
wire _00666_ ;
wire _00667_ ;
wire _00668_ ;
wire _00669_ ;
wire _00670_ ;
wire _00671_ ;
wire _00672_ ;
wire _00673_ ;
wire _00674_ ;
wire _00675_ ;
wire _00676_ ;
wire _00677_ ;
wire _00678_ ;
wire _00679_ ;
wire _00680_ ;
wire _00681_ ;
wire _00682_ ;
wire _00683_ ;
wire _00684_ ;
wire _00685_ ;
wire _00686_ ;
wire _00687_ ;
wire _00688_ ;
wire _00689_ ;
wire _00690_ ;
wire _00691_ ;
wire _00692_ ;
wire _00693_ ;
wire _00694_ ;
wire _00695_ ;
wire _00696_ ;
wire _00697_ ;
wire _00698_ ;
wire _00699_ ;
wire _00700_ ;
wire _00701_ ;
wire _00702_ ;
wire _00703_ ;
wire _00704_ ;
wire _00705_ ;
wire _00706_ ;
wire _00707_ ;
wire _00708_ ;
wire _00709_ ;
wire _00710_ ;
wire _00711_ ;
wire _00712_ ;
wire _00713_ ;
wire _00714_ ;
wire _00715_ ;
wire _00716_ ;
wire _00717_ ;
wire _00718_ ;
wire _00719_ ;
wire _00720_ ;
wire _00721_ ;
wire _00722_ ;
wire _00723_ ;
wire _00724_ ;
wire _00725_ ;
wire _00726_ ;
wire _00727_ ;
wire _00728_ ;
wire _00729_ ;
wire _00730_ ;
wire _00731_ ;
wire _00732_ ;
wire _00733_ ;
wire _00734_ ;
wire _00735_ ;
wire _00736_ ;
wire _00737_ ;
wire _00738_ ;
wire _00739_ ;
wire _00740_ ;
wire _00741_ ;
wire _00742_ ;
wire _00743_ ;
wire _00744_ ;
wire _00745_ ;
wire _00746_ ;
wire _00747_ ;
wire _00748_ ;
wire _00749_ ;
wire _00750_ ;
wire _00751_ ;
wire _00752_ ;
wire _00753_ ;
wire _00754_ ;
wire _00755_ ;
wire _00756_ ;
wire _00757_ ;
wire _00758_ ;
wire _00759_ ;
wire _00760_ ;
wire _00761_ ;
wire _00762_ ;
wire _00763_ ;
wire _00764_ ;
wire _00765_ ;
wire _00766_ ;
wire _00767_ ;
wire _00768_ ;
wire _00769_ ;
wire _00770_ ;
wire _00771_ ;
wire _00772_ ;
wire _00773_ ;
wire _00774_ ;
wire _00775_ ;
wire _00776_ ;
wire _00777_ ;
wire _00778_ ;
wire _00779_ ;
wire _00780_ ;
wire _00781_ ;
wire _00782_ ;
wire _00783_ ;
wire _00784_ ;
wire _00785_ ;
wire _00786_ ;
wire _00787_ ;
wire _00788_ ;
wire _00789_ ;
wire _00790_ ;
wire _00791_ ;
wire _00792_ ;
wire _00793_ ;
wire _00794_ ;
wire _00795_ ;
wire _00796_ ;
wire _00797_ ;
wire _00798_ ;
wire _00799_ ;
wire _00800_ ;
wire _00801_ ;
wire _00802_ ;
wire _00803_ ;
wire _00804_ ;
wire _00805_ ;
wire _00806_ ;
wire _00807_ ;
wire _00808_ ;
wire _00809_ ;
wire _00810_ ;
wire _00811_ ;
wire _00812_ ;
wire _00813_ ;
wire _00814_ ;
wire _00815_ ;
wire _00816_ ;
wire _00817_ ;
wire _00818_ ;
wire _00819_ ;
wire _00820_ ;
wire _00821_ ;
wire _00822_ ;
wire _00823_ ;
wire _00824_ ;
wire _00825_ ;
wire _00826_ ;
wire _00827_ ;
wire _00828_ ;
wire _00829_ ;
wire _00830_ ;
wire _00831_ ;
wire _00832_ ;
wire _00833_ ;
wire _00834_ ;
wire _00835_ ;
wire _00836_ ;
wire _00837_ ;
wire _00838_ ;
wire _00839_ ;
wire _00840_ ;
wire _00841_ ;
wire _00842_ ;
wire _00843_ ;
wire _00844_ ;
wire _00845_ ;
wire _00846_ ;
wire _00847_ ;
wire _00848_ ;
wire _00849_ ;
wire _00850_ ;
wire _00851_ ;
wire _00852_ ;
wire _00853_ ;
wire _00854_ ;
wire _00855_ ;
wire _00856_ ;
wire _00857_ ;
wire _00858_ ;
wire _00859_ ;
wire _00860_ ;
wire _00861_ ;
wire _00862_ ;
wire _00863_ ;
wire _00864_ ;
wire _00865_ ;
wire _00866_ ;
wire _00867_ ;
wire _00868_ ;
wire _00869_ ;
wire _00870_ ;
wire _00871_ ;
wire _00872_ ;
wire _00873_ ;
wire _00874_ ;
wire _00875_ ;
wire _00876_ ;
wire _00877_ ;
wire _00878_ ;
wire _00879_ ;
wire _00880_ ;
wire _00881_ ;
wire _00882_ ;
wire _00883_ ;
wire _00884_ ;
wire _00885_ ;
wire _00886_ ;
wire _00887_ ;
wire _00888_ ;
wire _00889_ ;
wire _00890_ ;
wire _00891_ ;
wire _00892_ ;
wire _00893_ ;
wire _00894_ ;
wire _00895_ ;
wire _00896_ ;
wire _00897_ ;
wire _00898_ ;
wire _00899_ ;
wire _00900_ ;
wire _00901_ ;
wire _00902_ ;
wire _00903_ ;
wire _00904_ ;
wire _00905_ ;
wire _00906_ ;
wire _00907_ ;
wire _00908_ ;
wire _00909_ ;
wire _00910_ ;
wire _00911_ ;
wire _00912_ ;
wire _00913_ ;
wire _00914_ ;
wire _00915_ ;
wire _00916_ ;
wire _00917_ ;
wire _00918_ ;
wire _00919_ ;
wire _00920_ ;
wire _00921_ ;
wire _00922_ ;
wire _00923_ ;
wire _00924_ ;
wire _00925_ ;
wire _00926_ ;
wire _00927_ ;
wire _00928_ ;
wire _00929_ ;
wire _00930_ ;
wire _00931_ ;
wire _00932_ ;
wire _00933_ ;
wire _00934_ ;
wire _00935_ ;
wire _00936_ ;
wire _00937_ ;
wire _00938_ ;
wire _00939_ ;
wire _00940_ ;
wire _00941_ ;
wire _00942_ ;
wire _00943_ ;
wire _00944_ ;
wire _00945_ ;
wire _00946_ ;
wire _00947_ ;
wire _00948_ ;
wire _00949_ ;
wire _00950_ ;
wire _00951_ ;
wire _00952_ ;
wire _00953_ ;
wire _00954_ ;
wire _00955_ ;
wire _00956_ ;
wire _00957_ ;
wire _00958_ ;
wire _00959_ ;
wire _00960_ ;
wire _00961_ ;
wire _00962_ ;
wire _00963_ ;
wire _00964_ ;
wire _00965_ ;
wire _00966_ ;
wire _00967_ ;
wire _00968_ ;
wire _00969_ ;
wire _00970_ ;
wire _00971_ ;
wire _00972_ ;
wire _00973_ ;
wire _00974_ ;
wire _00975_ ;
wire _00976_ ;
wire _00977_ ;
wire _00978_ ;
wire _00979_ ;
wire _00980_ ;
wire _00981_ ;
wire _00982_ ;
wire _00983_ ;
wire _00984_ ;
wire _00985_ ;
wire _00986_ ;
wire _00987_ ;
wire _00988_ ;
wire _00989_ ;
wire _00990_ ;
wire _00991_ ;
wire _00992_ ;
wire _00993_ ;
wire _00994_ ;
wire _00995_ ;
wire _00996_ ;
wire _00997_ ;
wire _00998_ ;
wire _00999_ ;
wire _01000_ ;
wire _01001_ ;
wire _01002_ ;
wire _01003_ ;
wire _01004_ ;
wire _01005_ ;
wire _01006_ ;
wire _01007_ ;
wire _01008_ ;
wire _01009_ ;
wire _01010_ ;
wire _01011_ ;
wire _01012_ ;
wire _01013_ ;
wire _01014_ ;
wire _01015_ ;
wire _01016_ ;
wire _01017_ ;
wire _01018_ ;
wire _01019_ ;
wire _01020_ ;
wire _01021_ ;
wire _01022_ ;
wire _01023_ ;
wire _01024_ ;
wire _01025_ ;
wire _01026_ ;
wire _01027_ ;
wire _01028_ ;
wire _01029_ ;
wire _01030_ ;
wire _01031_ ;
wire _01032_ ;
wire _01033_ ;
wire _01034_ ;
wire _01035_ ;
wire _01036_ ;
wire _01037_ ;
wire _01038_ ;
wire _01039_ ;
wire _01040_ ;
wire _01041_ ;
wire _01042_ ;
wire _01043_ ;
wire _01044_ ;
wire _01045_ ;
wire _01046_ ;
wire _01047_ ;
wire _01048_ ;
wire _01049_ ;
wire _01050_ ;
wire _01051_ ;
wire _01052_ ;
wire _01053_ ;
wire _01054_ ;
wire _01055_ ;
wire _01056_ ;
wire _01057_ ;
wire _01058_ ;
wire _01059_ ;
wire _01060_ ;
wire _01061_ ;
wire _01062_ ;
wire _01063_ ;
wire _01064_ ;
wire _01065_ ;
wire _01066_ ;
wire _01067_ ;
wire _01068_ ;
wire _01069_ ;
wire _01070_ ;
wire _01071_ ;
wire _01072_ ;
wire _01073_ ;
wire _01074_ ;
wire _01075_ ;
wire _01076_ ;
wire _01077_ ;
wire _01078_ ;
wire _01079_ ;
wire _01080_ ;
wire _01081_ ;
wire _01082_ ;
wire _01083_ ;
wire _01084_ ;
wire _01085_ ;
wire _01086_ ;
wire _01087_ ;
wire _01088_ ;
wire _01089_ ;
wire _01090_ ;
wire _01091_ ;
wire _01092_ ;
wire _01093_ ;
wire _01094_ ;
wire _01095_ ;
wire _01096_ ;
wire _01097_ ;
wire _01098_ ;
wire _01099_ ;
wire _01100_ ;
wire _01101_ ;
wire _01102_ ;
wire _01103_ ;
wire _01104_ ;
wire _01105_ ;
wire _01106_ ;
wire _01107_ ;
wire _01108_ ;
wire _01109_ ;
wire _01110_ ;
wire _01111_ ;
wire _01112_ ;
wire _01113_ ;
wire _01114_ ;
wire _01115_ ;
wire _01116_ ;
wire _01117_ ;
wire _01118_ ;
wire _01119_ ;
wire _01120_ ;
wire _01121_ ;
wire _01122_ ;
wire _01123_ ;
wire _01124_ ;
wire _01125_ ;
wire _01126_ ;
wire _01127_ ;
wire _01128_ ;
wire _01129_ ;
wire _01130_ ;
wire _01131_ ;
wire _01132_ ;
wire _01133_ ;
wire _01134_ ;
wire _01135_ ;
wire _01136_ ;
wire _01137_ ;
wire _01138_ ;
wire _01139_ ;
wire _01140_ ;
wire _01141_ ;
wire _01142_ ;
wire _01143_ ;
wire _01144_ ;
wire _01145_ ;
wire _01146_ ;
wire _01147_ ;
wire _01148_ ;
wire _01149_ ;
wire _01150_ ;
wire _01151_ ;
wire _01152_ ;
wire _01153_ ;
wire _01154_ ;
wire _01155_ ;
wire _01156_ ;
wire _01157_ ;
wire _01158_ ;
wire _01159_ ;
wire _01160_ ;
wire _01161_ ;
wire _01162_ ;
wire _01163_ ;
wire _01164_ ;
wire _01165_ ;
wire _01166_ ;
wire _01167_ ;
wire _01168_ ;
wire _01169_ ;
wire _01170_ ;
wire _01171_ ;
wire _01172_ ;
wire _01173_ ;
wire _01174_ ;
wire _01175_ ;
wire _01176_ ;
wire _01177_ ;
wire _01178_ ;
wire _01179_ ;
wire _01180_ ;
wire _01181_ ;
wire _01182_ ;
wire _01183_ ;
wire _01184_ ;
wire _01185_ ;
wire _01186_ ;
wire _01187_ ;
wire _01188_ ;
wire _01189_ ;
wire _01190_ ;
wire _01191_ ;
wire _01192_ ;
wire _01193_ ;
wire _01194_ ;
wire _01195_ ;
wire _01196_ ;
wire _01197_ ;
wire _01198_ ;
wire _01199_ ;
wire _01200_ ;
wire _01201_ ;
wire _01202_ ;
wire _01203_ ;
wire _01204_ ;
wire _01205_ ;
wire _01206_ ;
wire _01207_ ;
wire _01208_ ;
wire _01209_ ;
wire _01210_ ;
wire _01211_ ;
wire _01212_ ;
wire _01213_ ;
wire _01214_ ;
wire _01215_ ;
wire _01216_ ;
wire _01217_ ;
wire _01218_ ;
wire _01219_ ;
wire _01220_ ;
wire _01221_ ;
wire _01222_ ;
wire _01223_ ;
wire _01224_ ;
wire _01225_ ;
wire _01226_ ;
wire _01227_ ;
wire _01228_ ;
wire _01229_ ;
wire _01230_ ;
wire _01231_ ;
wire _01232_ ;
wire _01233_ ;
wire _01234_ ;
wire _01235_ ;
wire _01236_ ;
wire _01237_ ;
wire _01238_ ;
wire _01239_ ;
wire _01240_ ;
wire _01241_ ;
wire _01242_ ;
wire _01243_ ;
wire _01244_ ;
wire _01245_ ;
wire _01246_ ;
wire _01247_ ;
wire _01248_ ;
wire _01249_ ;
wire _01250_ ;
wire _01251_ ;
wire _01252_ ;
wire _01253_ ;
wire _01254_ ;
wire _01255_ ;
wire _01256_ ;
wire _01257_ ;
wire _01258_ ;
wire _01259_ ;
wire _01260_ ;
wire _01261_ ;
wire _01262_ ;
wire _01263_ ;
wire _01264_ ;
wire _01265_ ;
wire _01266_ ;
wire _01267_ ;
wire _01268_ ;
wire _01269_ ;
wire _01270_ ;
wire _01271_ ;
wire _01272_ ;
wire _01273_ ;
wire _01274_ ;
wire _01275_ ;
wire _01276_ ;
wire _01277_ ;
wire _01278_ ;
wire _01279_ ;
wire _01280_ ;
wire _01281_ ;
wire _01282_ ;
wire _01283_ ;
wire _01284_ ;
wire _01285_ ;
wire _01286_ ;
wire _01287_ ;
wire _01288_ ;
wire _01289_ ;
wire _01290_ ;
wire _01291_ ;
wire _01292_ ;
wire _01293_ ;
wire _01294_ ;
wire _01295_ ;
wire _01296_ ;
wire _01297_ ;
wire _01298_ ;
wire _01299_ ;
wire _01300_ ;
wire _01301_ ;
wire _01302_ ;
wire _01303_ ;
wire _01304_ ;
wire _01305_ ;
wire _01306_ ;
wire _01307_ ;
wire _01308_ ;
wire _01309_ ;
wire _01310_ ;
wire _01311_ ;
wire _01312_ ;
wire _01313_ ;
wire _01314_ ;
wire _01315_ ;
wire _01316_ ;
wire _01317_ ;
wire _01318_ ;
wire _01319_ ;
wire _01320_ ;
wire _01321_ ;
wire _01322_ ;
wire _01323_ ;
wire _01324_ ;
wire _01325_ ;
wire _01326_ ;
wire _01327_ ;
wire _01328_ ;
wire _01329_ ;
wire _01330_ ;
wire _01331_ ;
wire _01332_ ;
wire _01333_ ;
wire _01334_ ;
wire _01335_ ;
wire _01336_ ;
wire _01337_ ;
wire _01338_ ;
wire _01339_ ;
wire _01340_ ;
wire _01341_ ;
wire _01342_ ;
wire _01343_ ;
wire _01344_ ;
wire _01345_ ;
wire _01346_ ;
wire _01347_ ;
wire _01348_ ;
wire _01349_ ;
wire _01350_ ;
wire _01351_ ;
wire _01352_ ;
wire _01353_ ;
wire _01354_ ;
wire _01355_ ;
wire _01356_ ;
wire _01357_ ;
wire _01358_ ;
wire _01359_ ;
wire _01360_ ;
wire _01361_ ;
wire _01362_ ;
wire _01363_ ;
wire _01364_ ;
wire _01365_ ;
wire _01366_ ;
wire _01367_ ;
wire _01368_ ;
wire _01369_ ;
wire _01370_ ;
wire _01371_ ;
wire _01372_ ;
wire _01373_ ;
wire _01374_ ;
wire _01375_ ;
wire _01376_ ;
wire _01377_ ;
wire _01378_ ;
wire _01379_ ;
wire _01380_ ;
wire _01381_ ;
wire _01382_ ;
wire _01383_ ;
wire _01384_ ;
wire _01385_ ;
wire _01386_ ;
wire _01387_ ;
wire _01388_ ;
wire _01389_ ;
wire _01390_ ;
wire _01391_ ;
wire _01392_ ;
wire _01393_ ;
wire _01394_ ;
wire _01395_ ;
wire _01396_ ;
wire _01397_ ;
wire _01398_ ;
wire _01399_ ;
wire _01400_ ;
wire _01401_ ;
wire _01402_ ;
wire _01403_ ;
wire _01404_ ;
wire _01405_ ;
wire _01406_ ;
wire _01407_ ;
wire _01408_ ;
wire _01409_ ;
wire _01410_ ;
wire _01411_ ;
wire _01412_ ;
wire _01413_ ;
wire _01414_ ;
wire _01415_ ;
wire _01416_ ;
wire _01417_ ;
wire _01418_ ;
wire _01419_ ;
wire _01420_ ;
wire _01421_ ;
wire _01422_ ;
wire _01423_ ;
wire _01424_ ;
wire _01425_ ;
wire _01426_ ;
wire _01427_ ;
wire _01428_ ;
wire _01429_ ;
wire _01430_ ;
wire _01431_ ;
wire _01432_ ;
wire _01433_ ;
wire _01434_ ;
wire _01435_ ;
wire _01436_ ;
wire _01437_ ;
wire _01438_ ;
wire _01439_ ;
wire _01440_ ;
wire _01441_ ;
wire _01442_ ;
wire _01443_ ;
wire _01444_ ;
wire _01445_ ;
wire _01446_ ;
wire _01447_ ;
wire _01448_ ;
wire _01449_ ;
wire _01450_ ;
wire _01451_ ;
wire _01452_ ;
wire _01453_ ;
wire _01454_ ;
wire _01455_ ;
wire _01456_ ;
wire _01457_ ;
wire _01458_ ;
wire _01459_ ;
wire _01460_ ;
wire _01461_ ;
wire _01462_ ;
wire _01463_ ;
wire _01464_ ;
wire _01465_ ;
wire _01466_ ;
wire _01467_ ;
wire _01468_ ;
wire _01469_ ;
wire _01470_ ;
wire _01471_ ;
wire _01472_ ;
wire _01473_ ;
wire _01474_ ;
wire _01475_ ;
wire _01476_ ;
wire _01477_ ;
wire _01478_ ;
wire _01479_ ;
wire _01480_ ;
wire _01481_ ;
wire _01482_ ;
wire _01483_ ;
wire _01484_ ;
wire _01485_ ;
wire _01486_ ;
wire _01487_ ;
wire _01488_ ;
wire _01489_ ;
wire _01490_ ;
wire _01491_ ;
wire _01492_ ;
wire _01493_ ;
wire _01494_ ;
wire _01495_ ;
wire _01496_ ;
wire _01497_ ;
wire _01498_ ;
wire _01499_ ;
wire _01500_ ;
wire _01501_ ;
wire _01502_ ;
wire _01503_ ;
wire _01504_ ;
wire _01505_ ;
wire _01506_ ;
wire _01507_ ;
wire _01508_ ;
wire _01509_ ;
wire _01510_ ;
wire _01511_ ;
wire _01512_ ;
wire _01513_ ;
wire _01514_ ;
wire _01515_ ;
wire _01516_ ;
wire _01517_ ;
wire _01518_ ;
wire _01519_ ;
wire _01520_ ;
wire _01521_ ;
wire _01522_ ;
wire _01523_ ;
wire _01524_ ;
wire _01525_ ;
wire _01526_ ;
wire _01527_ ;
wire _01528_ ;
wire _01529_ ;
wire _01530_ ;
wire _01531_ ;
wire _01532_ ;
wire _01533_ ;
wire _01534_ ;
wire _01535_ ;
wire _01536_ ;
wire _01537_ ;
wire _01538_ ;
wire _01539_ ;
wire _01540_ ;
wire _01541_ ;
wire _01542_ ;
wire _01543_ ;
wire _01544_ ;
wire _01545_ ;
wire _01546_ ;
wire _01547_ ;
wire _01548_ ;
wire _01549_ ;
wire _01550_ ;
wire _01551_ ;
wire _01552_ ;
wire _01553_ ;
wire _01554_ ;
wire _01555_ ;
wire _01556_ ;
wire _01557_ ;
wire _01558_ ;
wire _01559_ ;
wire _01560_ ;
wire _01561_ ;
wire _01562_ ;
wire _01563_ ;
wire _01564_ ;
wire _01565_ ;
wire _01566_ ;
wire _01567_ ;
wire _01568_ ;
wire _01569_ ;
wire _01570_ ;
wire _01571_ ;
wire _01572_ ;
wire _01573_ ;
wire _01574_ ;
wire _01575_ ;
wire _01576_ ;
wire _01577_ ;
wire _01578_ ;
wire _01579_ ;
wire _01580_ ;
wire _01581_ ;
wire _01582_ ;
wire _01583_ ;
wire _01584_ ;
wire _01585_ ;
wire _01586_ ;
wire _01587_ ;
wire _01588_ ;
wire _01589_ ;
wire _01590_ ;
wire _01591_ ;
wire _01592_ ;
wire _01593_ ;
wire _01594_ ;
wire _01595_ ;
wire _01596_ ;
wire _01597_ ;
wire _01598_ ;
wire _01599_ ;
wire _01600_ ;
wire _01601_ ;
wire _01602_ ;
wire _01603_ ;
wire _01604_ ;
wire _01605_ ;
wire _01606_ ;
wire _01607_ ;
wire _01608_ ;
wire _01609_ ;
wire _01610_ ;
wire _01611_ ;
wire _01612_ ;
wire _01613_ ;
wire _01614_ ;
wire _01615_ ;
wire _01616_ ;
wire _01617_ ;
wire _01618_ ;
wire _01619_ ;
wire _01620_ ;
wire _01621_ ;
wire _01622_ ;
wire _01623_ ;
wire _01624_ ;
wire _01625_ ;
wire _01626_ ;
wire _01627_ ;
wire _01628_ ;
wire _01629_ ;
wire _01630_ ;
wire _01631_ ;
wire _01632_ ;
wire _01633_ ;
wire _01634_ ;
wire _01635_ ;
wire _01636_ ;
wire _01637_ ;
wire _01638_ ;
wire _01639_ ;
wire _01640_ ;
wire _01641_ ;
wire _01642_ ;
wire _01643_ ;
wire _01644_ ;
wire _01645_ ;
wire _01646_ ;
wire _01647_ ;
wire _01648_ ;
wire _01649_ ;
wire _01650_ ;
wire _01651_ ;
wire _01652_ ;
wire _01653_ ;
wire _01654_ ;
wire _01655_ ;
wire _01656_ ;
wire _01657_ ;
wire _01658_ ;
wire _01659_ ;
wire _01660_ ;
wire _01661_ ;
wire _01662_ ;
wire _01663_ ;
wire _01664_ ;
wire _01665_ ;
wire _01666_ ;
wire _01667_ ;
wire _01668_ ;
wire _01669_ ;
wire _01670_ ;
wire _01671_ ;
wire _01672_ ;
wire _01673_ ;
wire _01674_ ;
wire _01675_ ;
wire _01676_ ;
wire _01677_ ;
wire _01678_ ;
wire _01679_ ;
wire _01680_ ;
wire _01681_ ;
wire _01682_ ;
wire _01683_ ;
wire _01684_ ;
wire _01685_ ;
wire _01686_ ;
wire _01687_ ;
wire _01688_ ;
wire _01689_ ;
wire _01690_ ;
wire _01691_ ;
wire _01692_ ;
wire _01693_ ;
wire _01694_ ;
wire _01695_ ;
wire _01696_ ;
wire _01697_ ;
wire _01698_ ;
wire _01699_ ;
wire _01700_ ;
wire _01701_ ;
wire _01702_ ;
wire _01703_ ;
wire _01704_ ;
wire _01705_ ;
wire _01706_ ;
wire _01707_ ;
wire _01708_ ;
wire _01709_ ;
wire _01710_ ;
wire _01711_ ;
wire _01712_ ;
wire _01713_ ;
wire _01714_ ;
wire _01715_ ;
wire _01716_ ;
wire _01717_ ;
wire _01718_ ;
wire _01719_ ;
wire _01720_ ;
wire _01721_ ;
wire _01722_ ;
wire _01723_ ;
wire _01724_ ;
wire _01725_ ;
wire _01726_ ;
wire _01727_ ;
wire _01728_ ;
wire _01729_ ;
wire _01730_ ;
wire _01731_ ;
wire _01732_ ;
wire _01733_ ;
wire _01734_ ;
wire _01735_ ;
wire _01736_ ;
wire _01737_ ;
wire _01738_ ;
wire _01739_ ;
wire _01740_ ;
wire _01741_ ;
wire _01742_ ;
wire _01743_ ;
wire _01744_ ;
wire _01745_ ;
wire _01746_ ;
wire _01747_ ;
wire _01748_ ;
wire _01749_ ;
wire _01750_ ;
wire _01751_ ;
wire _01752_ ;
wire _01753_ ;
wire _01754_ ;
wire _01755_ ;
wire _01756_ ;
wire _01757_ ;
wire _01758_ ;
wire _01759_ ;
wire _01760_ ;
wire _01761_ ;
wire _01762_ ;
wire _01763_ ;
wire _01764_ ;
wire _01765_ ;
wire _01766_ ;
wire _01767_ ;
wire _01768_ ;
wire _01769_ ;
wire _01770_ ;
wire _01771_ ;
wire _01772_ ;
wire _01773_ ;
wire _01774_ ;
wire _01775_ ;
wire _01776_ ;
wire _01777_ ;
wire _01778_ ;
wire _01779_ ;
wire _01780_ ;
wire _01781_ ;
wire _01782_ ;
wire _01783_ ;
wire _01784_ ;
wire _01785_ ;
wire _01786_ ;
wire _01787_ ;
wire _01788_ ;
wire _01789_ ;
wire _01790_ ;
wire _01791_ ;
wire _01792_ ;
wire _01793_ ;
wire _01794_ ;
wire _01795_ ;
wire _01796_ ;
wire _01797_ ;
wire _01798_ ;
wire _01799_ ;
wire _01800_ ;
wire _01801_ ;
wire _01802_ ;
wire _01803_ ;
wire _01804_ ;
wire _01805_ ;
wire _01806_ ;
wire _01807_ ;
wire _01808_ ;
wire _01809_ ;
wire _01810_ ;
wire _01811_ ;
wire _01812_ ;
wire _01813_ ;
wire _01814_ ;
wire _01815_ ;
wire _01816_ ;
wire _01817_ ;
wire _01818_ ;
wire _01819_ ;
wire _01820_ ;
wire _01821_ ;
wire _01822_ ;
wire _01823_ ;
wire _01824_ ;
wire _01825_ ;
wire _01826_ ;
wire _01827_ ;
wire _01828_ ;
wire _01829_ ;
wire _01830_ ;
wire _01831_ ;
wire _01832_ ;
wire _01833_ ;
wire _01834_ ;
wire _01835_ ;
wire _01836_ ;
wire _01837_ ;
wire _01838_ ;
wire _01839_ ;
wire _01840_ ;
wire _01841_ ;
wire _01842_ ;
wire _01843_ ;
wire _01844_ ;
wire _01845_ ;
wire _01846_ ;
wire _01847_ ;
wire _01848_ ;
wire _01849_ ;
wire _01850_ ;
wire _01851_ ;
wire _01852_ ;
wire _01853_ ;
wire _01854_ ;
wire _01855_ ;
wire _01856_ ;
wire _01857_ ;
wire _01858_ ;
wire _01859_ ;
wire _01860_ ;
wire _01861_ ;
wire _01862_ ;
wire _01863_ ;
wire _01864_ ;
wire _01865_ ;
wire _01866_ ;
wire _01867_ ;
wire _01868_ ;
wire _01869_ ;
wire _01870_ ;
wire _01871_ ;
wire _01872_ ;
wire _01873_ ;
wire _01874_ ;
wire _01875_ ;
wire _01876_ ;
wire _01877_ ;
wire _01878_ ;
wire _01879_ ;
wire _01880_ ;
wire _01881_ ;
wire _01882_ ;
wire _01883_ ;
wire _01884_ ;
wire _01885_ ;
wire _01886_ ;
wire _01887_ ;
wire _01888_ ;
wire _01889_ ;
wire _01890_ ;
wire _01891_ ;
wire _01892_ ;
wire _01893_ ;
wire _01894_ ;
wire _01895_ ;
wire _01896_ ;
wire _01897_ ;
wire _01898_ ;
wire _01899_ ;
wire _01900_ ;
wire _01901_ ;
wire _01902_ ;
wire _01903_ ;
wire _01904_ ;
wire _01905_ ;
wire _01906_ ;
wire _01907_ ;
wire _01908_ ;
wire _01909_ ;
wire _01910_ ;
wire _01911_ ;
wire _01912_ ;
wire _01913_ ;
wire _01914_ ;
wire _01915_ ;
wire _01916_ ;
wire _01917_ ;
wire _01918_ ;
wire _01919_ ;
wire _01920_ ;
wire _01921_ ;
wire _01922_ ;
wire _01923_ ;
wire _01924_ ;
wire _01925_ ;
wire _01926_ ;
wire _01927_ ;
wire _01928_ ;
wire _01929_ ;
wire _01930_ ;
wire _01931_ ;
wire _01932_ ;
wire _01933_ ;
wire _01934_ ;
wire _01935_ ;
wire _01936_ ;
wire _01937_ ;
wire _01938_ ;
wire _01939_ ;
wire _01940_ ;
wire _01941_ ;
wire _01942_ ;
wire _01943_ ;
wire _01944_ ;
wire _01945_ ;
wire _01946_ ;
wire _01947_ ;
wire _01948_ ;
wire _01949_ ;
wire _01950_ ;
wire _01951_ ;
wire _01952_ ;
wire _01953_ ;
wire _01954_ ;
wire _01955_ ;
wire _01956_ ;
wire _01957_ ;
wire _01958_ ;
wire _01959_ ;
wire _01960_ ;
wire _01961_ ;
wire _01962_ ;
wire _01963_ ;
wire _01964_ ;
wire _01965_ ;
wire _01966_ ;
wire _01967_ ;
wire _01968_ ;
wire _01969_ ;
wire _01970_ ;
wire _01971_ ;
wire _01972_ ;
wire _01973_ ;
wire _01974_ ;
wire _01975_ ;
wire _01976_ ;
wire _01977_ ;
wire _01978_ ;
wire _01979_ ;
wire _01980_ ;
wire _01981_ ;
wire _01982_ ;
wire _01983_ ;
wire _01984_ ;
wire _01985_ ;
wire _01986_ ;
wire _01987_ ;
wire _01988_ ;
wire _01989_ ;
wire _01990_ ;
wire _01991_ ;
wire _01992_ ;
wire _01993_ ;
wire _01994_ ;
wire _01995_ ;
wire _01996_ ;
wire _01997_ ;
wire _01998_ ;
wire _01999_ ;
wire _02000_ ;
wire _02001_ ;
wire _02002_ ;
wire _02003_ ;
wire _02004_ ;
wire _02005_ ;
wire _02006_ ;
wire _02007_ ;
wire _02008_ ;
wire _02009_ ;
wire _02010_ ;
wire _02011_ ;
wire _02012_ ;
wire _02013_ ;
wire _02014_ ;
wire _02015_ ;
wire _02016_ ;
wire _02017_ ;
wire _02018_ ;
wire _02019_ ;
wire _02020_ ;
wire _02021_ ;
wire _02022_ ;
wire _02023_ ;
wire _02024_ ;
wire _02025_ ;
wire _02026_ ;
wire _02027_ ;
wire _02028_ ;
wire _02029_ ;
wire _02030_ ;
wire _02031_ ;
wire _02032_ ;
wire _02033_ ;
wire _02034_ ;
wire _02035_ ;
wire _02036_ ;
wire _02037_ ;
wire _02038_ ;
wire _02039_ ;
wire _02040_ ;
wire _02041_ ;
wire _02042_ ;
wire _02043_ ;
wire _02044_ ;
wire _02045_ ;
wire _02046_ ;
wire _02047_ ;
wire _02048_ ;
wire _02049_ ;
wire _02050_ ;
wire _02051_ ;
wire _02052_ ;
wire _02053_ ;
wire _02054_ ;
wire _02055_ ;
wire _02056_ ;
wire _02057_ ;
wire _02058_ ;
wire _02059_ ;
wire _02060_ ;
wire _02061_ ;
wire _02062_ ;
wire _02063_ ;
wire _02064_ ;
wire _02065_ ;
wire _02066_ ;
wire _02067_ ;
wire _02068_ ;
wire _02069_ ;
wire _02070_ ;
wire _02071_ ;
wire _02072_ ;
wire _02073_ ;
wire _02074_ ;
wire _02075_ ;
wire _02076_ ;
wire _02077_ ;
wire _02078_ ;
wire _02079_ ;
wire _02080_ ;
wire _02081_ ;
wire _02082_ ;
wire _02083_ ;
wire _02084_ ;
wire _02085_ ;
wire _02086_ ;
wire _02087_ ;
wire _02088_ ;
wire _02089_ ;
wire _02090_ ;
wire _02091_ ;
wire _02092_ ;
wire _02093_ ;
wire _02094_ ;
wire _02095_ ;
wire _02096_ ;
wire _02097_ ;
wire _02098_ ;
wire _02099_ ;
wire _02100_ ;
wire _02101_ ;
wire _02102_ ;
wire _02103_ ;
wire _02104_ ;
wire _02105_ ;
wire _02106_ ;
wire _02107_ ;
wire _02108_ ;
wire _02109_ ;
wire _02110_ ;
wire _02111_ ;
wire _02112_ ;
wire _02113_ ;
wire _02114_ ;
wire _02115_ ;
wire _02116_ ;
wire _02117_ ;
wire _02118_ ;
wire _02119_ ;
wire _02120_ ;
wire _02121_ ;
wire _02122_ ;
wire _02123_ ;
wire _02124_ ;
wire _02125_ ;
wire _02126_ ;
wire _02127_ ;
wire _02128_ ;
wire _02129_ ;
wire _02130_ ;
wire _02131_ ;
wire _02132_ ;
wire _02133_ ;
wire _02134_ ;
wire _02135_ ;
wire _02136_ ;
wire _02137_ ;
wire _02138_ ;
wire _02139_ ;
wire _02140_ ;
wire _02141_ ;
wire _02142_ ;
wire _02143_ ;
wire _02144_ ;
wire _02145_ ;
wire _02146_ ;
wire _02147_ ;
wire _02148_ ;
wire _02149_ ;
wire _02150_ ;
wire _02151_ ;
wire _02152_ ;
wire _02153_ ;
wire _02154_ ;
wire _02155_ ;
wire _02156_ ;
wire _02157_ ;
wire _02158_ ;
wire _02159_ ;
wire _02160_ ;
wire _02161_ ;
wire _02162_ ;
wire _02163_ ;
wire _02164_ ;
wire _02165_ ;
wire _02166_ ;
wire _02167_ ;
wire _02168_ ;
wire _02169_ ;
wire _02170_ ;
wire _02171_ ;
wire _02172_ ;
wire _02173_ ;
wire _02174_ ;
wire _02175_ ;
wire _02176_ ;
wire _02177_ ;
wire _02178_ ;
wire _02179_ ;
wire _02180_ ;
wire _02181_ ;
wire _02182_ ;
wire _02183_ ;
wire _02184_ ;
wire _02185_ ;
wire _02186_ ;
wire _02187_ ;
wire _02188_ ;
wire _02189_ ;
wire _02190_ ;
wire _02191_ ;
wire _02192_ ;
wire _02193_ ;
wire _02194_ ;
wire _02195_ ;
wire _02196_ ;
wire _02197_ ;
wire _02198_ ;
wire _02199_ ;
wire _02200_ ;
wire _02201_ ;
wire _02202_ ;
wire _02203_ ;
wire _02204_ ;
wire _02205_ ;
wire _02206_ ;
wire _02207_ ;
wire _02208_ ;
wire _02209_ ;
wire _02210_ ;
wire _02211_ ;
wire _02212_ ;
wire _02213_ ;
wire _02214_ ;
wire _02215_ ;
wire _02216_ ;
wire _02217_ ;
wire _02218_ ;
wire _02219_ ;
wire _02220_ ;
wire _02221_ ;
wire _02222_ ;
wire _02223_ ;
wire _02224_ ;
wire _02225_ ;
wire _02226_ ;
wire _02227_ ;
wire _02228_ ;
wire _02229_ ;
wire _02230_ ;
wire _02231_ ;
wire _02232_ ;
wire _02233_ ;
wire _02234_ ;
wire _02235_ ;
wire _02236_ ;
wire _02237_ ;
wire _02238_ ;
wire _02239_ ;
wire _02240_ ;
wire _02241_ ;
wire _02242_ ;
wire _02243_ ;
wire _02244_ ;
wire _02245_ ;
wire _02246_ ;
wire _02247_ ;
wire _02248_ ;
wire _02249_ ;
wire _02250_ ;
wire _02251_ ;
wire _02252_ ;
wire _02253_ ;
wire _02254_ ;
wire _02255_ ;
wire _02256_ ;
wire _02257_ ;
wire _02258_ ;
wire _02259_ ;
wire _02260_ ;
wire _02261_ ;
wire _02262_ ;
wire _02263_ ;
wire _02264_ ;
wire _02265_ ;
wire _02266_ ;
wire _02267_ ;
wire _02268_ ;
wire _02269_ ;
wire _02270_ ;
wire _02271_ ;
wire _02272_ ;
wire _02273_ ;
wire _02274_ ;
wire _02275_ ;
wire _02276_ ;
wire _02277_ ;
wire _02278_ ;
wire _02279_ ;
wire _02280_ ;
wire _02281_ ;
wire _02282_ ;
wire _02283_ ;
wire _02284_ ;
wire _02285_ ;
wire _02286_ ;
wire _02287_ ;
wire _02288_ ;
wire _02289_ ;
wire _02290_ ;
wire _02291_ ;
wire _02292_ ;
wire _02293_ ;
wire _02294_ ;
wire _02295_ ;
wire _02296_ ;
wire _02297_ ;
wire _02298_ ;
wire _02299_ ;
wire _02300_ ;
wire _02301_ ;
wire _02302_ ;
wire _02303_ ;
wire _02304_ ;
wire _02305_ ;
wire _02306_ ;
wire _02307_ ;
wire _02308_ ;
wire _02309_ ;
wire _02310_ ;
wire _02311_ ;
wire _02312_ ;
wire _02313_ ;
wire _02314_ ;
wire _02315_ ;
wire _02316_ ;
wire _02317_ ;
wire _02318_ ;
wire _02319_ ;
wire _02320_ ;
wire _02321_ ;
wire _02322_ ;
wire _02323_ ;
wire _02324_ ;
wire _02325_ ;
wire _02326_ ;
wire _02327_ ;
wire _02328_ ;
wire _02329_ ;
wire _02330_ ;
wire _02331_ ;
wire _02332_ ;
wire _02333_ ;
wire _02334_ ;
wire _02335_ ;
wire _02336_ ;
wire _02337_ ;
wire _02338_ ;
wire _02339_ ;
wire _02340_ ;
wire _02341_ ;
wire _02342_ ;
wire _02343_ ;
wire _02344_ ;
wire _02345_ ;
wire _02346_ ;
wire _02347_ ;
wire _02348_ ;
wire _02349_ ;
wire _02350_ ;
wire _02351_ ;
wire _02352_ ;
wire _02353_ ;
wire _02354_ ;
wire _02355_ ;
wire _02356_ ;
wire _02357_ ;
wire _02358_ ;
wire _02359_ ;
wire _02360_ ;
wire _02361_ ;
wire _02362_ ;
wire _02363_ ;
wire _02364_ ;
wire _02365_ ;
wire _02366_ ;
wire _02367_ ;
wire _02368_ ;
wire _02369_ ;
wire _02370_ ;
wire _02371_ ;
wire _02372_ ;
wire _02373_ ;
wire _02374_ ;
wire _02375_ ;
wire _02376_ ;
wire _02377_ ;
wire _02378_ ;
wire _02379_ ;
wire _02380_ ;
wire _02381_ ;
wire _02382_ ;
wire _02383_ ;
wire _02384_ ;
wire _02385_ ;
wire _02386_ ;
wire _02387_ ;
wire _02388_ ;
wire _02389_ ;
wire _02390_ ;
wire _02391_ ;
wire _02392_ ;
wire _02393_ ;
wire _02394_ ;
wire _02395_ ;
wire _02396_ ;
wire _02397_ ;
wire _02398_ ;
wire _02399_ ;
wire _02400_ ;
wire _02401_ ;
wire _02402_ ;
wire _02403_ ;
wire _02404_ ;
wire _02405_ ;
wire _02406_ ;
wire _02407_ ;
wire _02408_ ;
wire _02409_ ;
wire _02410_ ;
wire _02411_ ;
wire _02412_ ;
wire _02413_ ;
wire _02414_ ;
wire _02415_ ;
wire _02416_ ;
wire _02417_ ;
wire _02418_ ;
wire _02419_ ;
wire _02420_ ;
wire _02421_ ;
wire _02422_ ;
wire _02423_ ;
wire _02424_ ;
wire _02425_ ;
wire _02426_ ;
wire _02427_ ;
wire _02428_ ;
wire _02429_ ;
wire _02430_ ;
wire _02431_ ;
wire _02432_ ;
wire _02433_ ;
wire _02434_ ;
wire _02435_ ;
wire _02436_ ;
wire _02437_ ;
wire _02438_ ;
wire _02439_ ;
wire _02440_ ;
wire _02441_ ;
wire _02442_ ;
wire _02443_ ;
wire _02444_ ;
wire _02445_ ;
wire _02446_ ;
wire _02447_ ;
wire _02448_ ;
wire _02449_ ;
wire _02450_ ;
wire _02451_ ;
wire _02452_ ;
wire _02453_ ;
wire _02454_ ;
wire _02455_ ;
wire _02456_ ;
wire _02457_ ;
wire _02458_ ;
wire _02459_ ;
wire _02460_ ;
wire _02461_ ;
wire _02462_ ;
wire _02463_ ;
wire _02464_ ;
wire _02465_ ;
wire _02466_ ;
wire _02467_ ;
wire _02468_ ;
wire _02469_ ;
wire _02470_ ;
wire _02471_ ;
wire _02472_ ;
wire _02473_ ;
wire _02474_ ;
wire _02475_ ;
wire _02476_ ;
wire _02477_ ;
wire _02478_ ;
wire _02479_ ;
wire _02480_ ;
wire _02481_ ;
wire _02482_ ;
wire _02483_ ;
wire _02484_ ;
wire _02485_ ;
wire _02486_ ;
wire _02487_ ;
wire _02488_ ;
wire _02489_ ;
wire _02490_ ;
wire _02491_ ;
wire _02492_ ;
wire _02493_ ;
wire _02494_ ;
wire _02495_ ;
wire _02496_ ;
wire _02497_ ;
wire _02498_ ;
wire _02499_ ;
wire _02500_ ;
wire _02501_ ;
wire _02502_ ;
wire _02503_ ;
wire _02504_ ;
wire _02505_ ;
wire _02506_ ;
wire _02507_ ;
wire _02508_ ;
wire _02509_ ;
wire _02510_ ;
wire _02511_ ;
wire _02512_ ;
wire _02513_ ;
wire _02514_ ;
wire _02515_ ;
wire _02516_ ;
wire _02517_ ;
wire _02518_ ;
wire _02519_ ;
wire _02520_ ;
wire _02521_ ;
wire _02522_ ;
wire _02523_ ;
wire _02524_ ;
wire _02525_ ;
wire _02526_ ;
wire _02527_ ;
wire _02528_ ;
wire _02529_ ;
wire _02530_ ;
wire _02531_ ;
wire _02532_ ;
wire _02533_ ;
wire _02534_ ;
wire _02535_ ;
wire _02536_ ;
wire _02537_ ;
wire _02538_ ;
wire _02539_ ;
wire _02540_ ;
wire _02541_ ;
wire _02542_ ;
wire _02543_ ;
wire _02544_ ;
wire _02545_ ;
wire _02546_ ;
wire _02547_ ;
wire _02548_ ;
wire _02549_ ;
wire _02550_ ;
wire _02551_ ;
wire _02552_ ;
wire _02553_ ;
wire _02554_ ;
wire _02555_ ;
wire _02556_ ;
wire _02557_ ;
wire _02558_ ;
wire _02559_ ;
wire _02560_ ;
wire _02561_ ;
wire _02562_ ;
wire _02563_ ;
wire _02564_ ;
wire _02565_ ;
wire _02566_ ;
wire _02567_ ;
wire _02568_ ;
wire _02569_ ;
wire _02570_ ;
wire _02571_ ;
wire _02572_ ;
wire _02573_ ;
wire _02574_ ;
wire _02575_ ;
wire _02576_ ;
wire _02577_ ;
wire _02578_ ;
wire _02579_ ;
wire _02580_ ;
wire _02581_ ;
wire _02582_ ;
wire _02583_ ;
wire _02584_ ;
wire _02585_ ;
wire _02586_ ;
wire _02587_ ;
wire _02588_ ;
wire _02589_ ;
wire _02590_ ;
wire _02591_ ;
wire _02592_ ;
wire _02593_ ;
wire _02594_ ;
wire _02595_ ;
wire _02596_ ;
wire _02597_ ;
wire _02598_ ;
wire _02599_ ;
wire _02600_ ;
wire _02601_ ;
wire _02602_ ;
wire _02603_ ;
wire _02604_ ;
wire _02605_ ;
wire _02606_ ;
wire _02607_ ;
wire _02608_ ;
wire _02609_ ;
wire _02610_ ;
wire _02611_ ;
wire _02612_ ;
wire _02613_ ;
wire _02614_ ;
wire _02615_ ;
wire _02616_ ;
wire _02617_ ;
wire _02618_ ;
wire _02619_ ;
wire _02620_ ;
wire _02621_ ;
wire _02622_ ;
wire _02623_ ;
wire _02624_ ;
wire _02625_ ;
wire _02626_ ;
wire _02627_ ;
wire _02628_ ;
wire _02629_ ;
wire _02630_ ;
wire _02631_ ;
wire _02632_ ;
wire _02633_ ;
wire _02634_ ;
wire _02635_ ;
wire _02636_ ;
wire _02637_ ;
wire _02638_ ;
wire _02639_ ;
wire _02640_ ;
wire _02641_ ;
wire _02642_ ;
wire _02643_ ;
wire _02644_ ;
wire _02645_ ;
wire _02646_ ;
wire _02647_ ;
wire _02648_ ;
wire _02649_ ;
wire _02650_ ;
wire _02651_ ;
wire _02652_ ;
wire _02653_ ;
wire _02654_ ;
wire _02655_ ;
wire _02656_ ;
wire _02657_ ;
wire _02658_ ;
wire _02659_ ;
wire _02660_ ;
wire _02661_ ;
wire _02662_ ;
wire _02663_ ;
wire _02664_ ;
wire _02665_ ;
wire _02666_ ;
wire _02667_ ;
wire _02668_ ;
wire _02669_ ;
wire _02670_ ;
wire _02671_ ;
wire _02672_ ;
wire _02673_ ;
wire _02674_ ;
wire _02675_ ;
wire _02676_ ;
wire _02677_ ;
wire _02678_ ;
wire _02679_ ;
wire _02680_ ;
wire _02681_ ;
wire _02682_ ;
wire _02683_ ;
wire _02684_ ;
wire _02685_ ;
wire _02686_ ;
wire _02687_ ;
wire _02688_ ;
wire _02689_ ;
wire _02690_ ;
wire _02691_ ;
wire _02692_ ;
wire _02693_ ;
wire _02694_ ;
wire _02695_ ;
wire _02696_ ;
wire _02697_ ;
wire _02698_ ;
wire _02699_ ;
wire _02700_ ;
wire _02701_ ;
wire _02702_ ;
wire _02703_ ;
wire _02704_ ;
wire _02705_ ;
wire _02706_ ;
wire _02707_ ;
wire _02708_ ;
wire _02709_ ;
wire _02710_ ;
wire _02711_ ;
wire _02712_ ;
wire _02713_ ;
wire _02714_ ;
wire _02715_ ;
wire _02716_ ;
wire _02717_ ;
wire _02718_ ;
wire _02719_ ;
wire _02720_ ;
wire _02721_ ;
wire _02722_ ;
wire _02723_ ;
wire _02724_ ;
wire _02725_ ;
wire _02726_ ;
wire _02727_ ;
wire _02728_ ;
wire _02729_ ;
wire _02730_ ;
wire _02731_ ;
wire _02732_ ;
wire _02733_ ;
wire _02734_ ;
wire _02735_ ;
wire _02736_ ;
wire _02737_ ;
wire _02738_ ;
wire _02739_ ;
wire _02740_ ;
wire _02741_ ;
wire _02742_ ;
wire _02743_ ;
wire _02744_ ;
wire _02745_ ;
wire _02746_ ;
wire _02747_ ;
wire _02748_ ;
wire _02749_ ;
wire _02750_ ;
wire _02751_ ;
wire _02752_ ;
wire _02753_ ;
wire _02754_ ;
wire _02755_ ;
wire _02756_ ;
wire _02757_ ;
wire _02758_ ;
wire _02759_ ;
wire _02760_ ;
wire _02761_ ;
wire _02762_ ;
wire _02763_ ;
wire _02764_ ;
wire _02765_ ;
wire _02766_ ;
wire _02767_ ;
wire _02768_ ;
wire _02769_ ;
wire _02770_ ;
wire _02771_ ;
wire _02772_ ;
wire _02773_ ;
wire _02774_ ;
wire _02775_ ;
wire _02776_ ;
wire _02777_ ;
wire _02778_ ;
wire _02779_ ;
wire _02780_ ;
wire _02781_ ;
wire _02782_ ;
wire _02783_ ;
wire _02784_ ;
wire _02785_ ;
wire _02786_ ;
wire _02787_ ;
wire _02788_ ;
wire _02789_ ;
wire _02790_ ;
wire _02791_ ;
wire _02792_ ;
wire _02793_ ;
wire _02794_ ;
wire _02795_ ;
wire _02796_ ;
wire _02797_ ;
wire _02798_ ;
wire _02799_ ;
wire _02800_ ;
wire _02801_ ;
wire _02802_ ;
wire _02803_ ;
wire _02804_ ;
wire _02805_ ;
wire _02806_ ;
wire _02807_ ;
wire _02808_ ;
wire _02809_ ;
wire _02810_ ;
wire _02811_ ;
wire _02812_ ;
wire _02813_ ;
wire _02814_ ;
wire _02815_ ;
wire _02816_ ;
wire _02817_ ;
wire _02818_ ;
wire _02819_ ;
wire _02820_ ;
wire _02821_ ;
wire _02822_ ;
wire _02823_ ;
wire _02824_ ;
wire _02825_ ;
wire _02826_ ;
wire _02827_ ;
wire _02828_ ;
wire _02829_ ;
wire _02830_ ;
wire _02831_ ;
wire _02832_ ;
wire _02833_ ;
wire _02834_ ;
wire _02835_ ;
wire _02836_ ;
wire _02837_ ;
wire _02838_ ;
wire _02839_ ;
wire _02840_ ;
wire _02841_ ;
wire _02842_ ;
wire _02843_ ;
wire _02844_ ;
wire _02845_ ;
wire _02846_ ;
wire _02847_ ;
wire _02848_ ;
wire _02849_ ;
wire _02850_ ;
wire _02851_ ;
wire _02852_ ;
wire _02853_ ;
wire _02854_ ;
wire _02855_ ;
wire _02856_ ;
wire _02857_ ;
wire _02858_ ;
wire _02859_ ;
wire _02860_ ;
wire _02861_ ;
wire _02862_ ;
wire _02863_ ;
wire _02864_ ;
wire _02865_ ;
wire _02866_ ;
wire _02867_ ;
wire _02868_ ;
wire _02869_ ;
wire _02870_ ;
wire _02871_ ;
wire _02872_ ;
wire _02873_ ;
wire _02874_ ;
wire _02875_ ;
wire _02876_ ;
wire _02877_ ;
wire _02878_ ;
wire _02879_ ;
wire _02880_ ;
wire _02881_ ;
wire _02882_ ;
wire _02883_ ;
wire _02884_ ;
wire _02885_ ;
wire _02886_ ;
wire _02887_ ;
wire _02888_ ;
wire _02889_ ;
wire _02890_ ;
wire _02891_ ;
wire _02892_ ;
wire _02893_ ;
wire _02894_ ;
wire _02895_ ;
wire _02896_ ;
wire _02897_ ;
wire _02898_ ;
wire _02899_ ;
wire _02900_ ;
wire _02901_ ;
wire _02902_ ;
wire _02903_ ;
wire _02904_ ;
wire _02905_ ;
wire _02906_ ;
wire _02907_ ;
wire _02908_ ;
wire _02909_ ;
wire _02910_ ;
wire _02911_ ;
wire _02912_ ;
wire _02913_ ;
wire _02914_ ;
wire _02915_ ;
wire _02916_ ;
wire _02917_ ;
wire _02918_ ;
wire _02919_ ;
wire _02920_ ;
wire _02921_ ;
wire _02922_ ;
wire _02923_ ;
wire _02924_ ;
wire _02925_ ;
wire _02926_ ;
wire _02927_ ;
wire _02928_ ;
wire _02929_ ;
wire _02930_ ;
wire _02931_ ;
wire _02932_ ;
wire _02933_ ;
wire _02934_ ;
wire _02935_ ;
wire _02936_ ;
wire _02937_ ;
wire _02938_ ;
wire _02939_ ;
wire _02940_ ;
wire _02941_ ;
wire _02942_ ;
wire _02943_ ;
wire _02944_ ;
wire _02945_ ;
wire _02946_ ;
wire _02947_ ;
wire _02948_ ;
wire _02949_ ;
wire _02950_ ;
wire _02951_ ;
wire _02952_ ;
wire _02953_ ;
wire _02954_ ;
wire _02955_ ;
wire _02956_ ;
wire _02957_ ;
wire _02958_ ;
wire _02959_ ;
wire _02960_ ;
wire _02961_ ;
wire _02962_ ;
wire _02963_ ;
wire _02964_ ;
wire _02965_ ;
wire _02966_ ;
wire _02967_ ;
wire _02968_ ;
wire _02969_ ;
wire _02970_ ;
wire _02971_ ;
wire _02972_ ;
wire _02973_ ;
wire _02974_ ;
wire _02975_ ;
wire _02976_ ;
wire _02977_ ;
wire _02978_ ;
wire _02979_ ;
wire _02980_ ;
wire _02981_ ;
wire _02982_ ;
wire _02983_ ;
wire _02984_ ;
wire _02985_ ;
wire _02986_ ;
wire _02987_ ;
wire _02988_ ;
wire _02989_ ;
wire _02990_ ;
wire _02991_ ;
wire _02992_ ;
wire _02993_ ;
wire _02994_ ;
wire _02995_ ;
wire _02996_ ;
wire _02997_ ;
wire _02998_ ;
wire _02999_ ;
wire _03000_ ;
wire _03001_ ;
wire _03002_ ;
wire _03003_ ;
wire _03004_ ;
wire _03005_ ;
wire _03006_ ;
wire _03007_ ;
wire _03008_ ;
wire _03009_ ;
wire _03010_ ;
wire _03011_ ;
wire _03012_ ;
wire _03013_ ;
wire _03014_ ;
wire _03015_ ;
wire _03016_ ;
wire _03017_ ;
wire _03018_ ;
wire _03019_ ;
wire _03020_ ;
wire _03021_ ;
wire _03022_ ;
wire _03023_ ;
wire _03024_ ;
wire _03025_ ;
wire _03026_ ;
wire _03027_ ;
wire _03028_ ;
wire _03029_ ;
wire _03030_ ;
wire _03031_ ;
wire _03032_ ;
wire _03033_ ;
wire _03034_ ;
wire _03035_ ;
wire _03036_ ;
wire _03037_ ;
wire _03038_ ;
wire _03039_ ;
wire _03040_ ;
wire _03041_ ;
wire _03042_ ;
wire _03043_ ;
wire _03044_ ;
wire _03045_ ;
wire _03046_ ;
wire _03047_ ;
wire _03048_ ;
wire _03049_ ;
wire _03050_ ;
wire _03051_ ;
wire _03052_ ;
wire _03053_ ;
wire _03054_ ;
wire _03055_ ;
wire _03056_ ;
wire _03057_ ;
wire _03058_ ;
wire _03059_ ;
wire _03060_ ;
wire _03061_ ;
wire _03062_ ;
wire _03063_ ;
wire _03064_ ;
wire _03065_ ;
wire _03066_ ;
wire _03067_ ;
wire _03068_ ;
wire _03069_ ;
wire _03070_ ;
wire _03071_ ;
wire _03072_ ;
wire _03073_ ;
wire _03074_ ;
wire _03075_ ;
wire _03076_ ;
wire _03077_ ;
wire _03078_ ;
wire _03079_ ;
wire _03080_ ;
wire _03081_ ;
wire _03082_ ;
wire _03083_ ;
wire _03084_ ;
wire _03085_ ;
wire _03086_ ;
wire _03087_ ;
wire _03088_ ;
wire _03089_ ;
wire _03090_ ;
wire _03091_ ;
wire _03092_ ;
wire _03093_ ;
wire _03094_ ;
wire _03095_ ;
wire _03096_ ;
wire _03097_ ;
wire _03098_ ;
wire _03099_ ;
wire _03100_ ;
wire _03101_ ;
wire _03102_ ;
wire _03103_ ;
wire _03104_ ;
wire _03105_ ;
wire _03106_ ;
wire _03107_ ;
wire _03108_ ;
wire _03109_ ;
wire _03110_ ;
wire _03111_ ;
wire _03112_ ;
wire _03113_ ;
wire _03114_ ;
wire _03115_ ;
wire _03116_ ;
wire _03117_ ;
wire _03118_ ;
wire _03119_ ;
wire _03120_ ;
wire _03121_ ;
wire _03122_ ;
wire _03123_ ;
wire _03124_ ;
wire _03125_ ;
wire _03126_ ;
wire _03127_ ;
wire _03128_ ;
wire _03129_ ;
wire _03130_ ;
wire _03131_ ;
wire _03132_ ;
wire _03133_ ;
wire _03134_ ;
wire _03135_ ;
wire _03136_ ;
wire _03137_ ;
wire _03138_ ;
wire _03139_ ;
wire _03140_ ;
wire _03141_ ;
wire _03142_ ;
wire _03143_ ;
wire _03144_ ;
wire _03145_ ;
wire _03146_ ;
wire _03147_ ;
wire _03148_ ;
wire _03149_ ;
wire _03150_ ;
wire _03151_ ;
wire _03152_ ;
wire _03153_ ;
wire _03154_ ;
wire _03155_ ;
wire _03156_ ;
wire _03157_ ;
wire _03158_ ;
wire _03159_ ;
wire _03160_ ;
wire _03161_ ;
wire _03162_ ;
wire _03163_ ;
wire _03164_ ;
wire _03165_ ;
wire _03166_ ;
wire _03167_ ;
wire _03168_ ;
wire _03169_ ;
wire _03170_ ;
wire _03171_ ;
wire _03172_ ;
wire _03173_ ;
wire _03174_ ;
wire _03175_ ;
wire _03176_ ;
wire _03177_ ;
wire _03178_ ;
wire _03179_ ;
wire _03180_ ;
wire _03181_ ;
wire _03182_ ;
wire _03183_ ;
wire _03184_ ;
wire _03185_ ;
wire _03186_ ;
wire _03187_ ;
wire _03188_ ;
wire _03189_ ;
wire _03190_ ;
wire _03191_ ;
wire _03192_ ;
wire _03193_ ;
wire _03194_ ;
wire _03195_ ;
wire _03196_ ;
wire _03197_ ;
wire _03198_ ;
wire _03199_ ;
wire _03200_ ;
wire _03201_ ;
wire _03202_ ;
wire _03203_ ;
wire _03204_ ;
wire _03205_ ;
wire _03206_ ;
wire _03207_ ;
wire _03208_ ;
wire _03209_ ;
wire _03210_ ;
wire _03211_ ;
wire _03212_ ;
wire _03213_ ;
wire _03214_ ;
wire _03215_ ;
wire _03216_ ;
wire _03217_ ;
wire _03218_ ;
wire _03219_ ;
wire _03220_ ;
wire _03221_ ;
wire _03222_ ;
wire _03223_ ;
wire _03224_ ;
wire _03225_ ;
wire _03226_ ;
wire _03227_ ;
wire _03228_ ;
wire _03229_ ;
wire _03230_ ;
wire _03231_ ;
wire _03232_ ;
wire _03233_ ;
wire _03234_ ;
wire _03235_ ;
wire _03236_ ;
wire _03237_ ;
wire _03238_ ;
wire _03239_ ;
wire _03240_ ;
wire _03241_ ;
wire _03242_ ;
wire _03243_ ;
wire _03244_ ;
wire _03245_ ;
wire _03246_ ;
wire _03247_ ;
wire _03248_ ;
wire _03249_ ;
wire _03250_ ;
wire _03251_ ;
wire _03252_ ;
wire _03253_ ;
wire _03254_ ;
wire _03255_ ;
wire _03256_ ;
wire _03257_ ;
wire _03258_ ;
wire _03259_ ;
wire _03260_ ;
wire _03261_ ;
wire _03262_ ;
wire _03263_ ;
wire _03264_ ;
wire _03265_ ;
wire _03266_ ;
wire _03267_ ;
wire _03268_ ;
wire _03269_ ;
wire _03270_ ;
wire _03271_ ;
wire _03272_ ;
wire _03273_ ;
wire _03274_ ;
wire _03275_ ;
wire _03276_ ;
wire _03277_ ;
wire _03278_ ;
wire _03279_ ;
wire _03280_ ;
wire _03281_ ;
wire _03282_ ;
wire _03283_ ;
wire _03284_ ;
wire _03285_ ;
wire _03286_ ;
wire _03287_ ;
wire _03288_ ;
wire _03289_ ;
wire _03290_ ;
wire _03291_ ;
wire _03292_ ;
wire _03293_ ;
wire _03294_ ;
wire _03295_ ;
wire _03296_ ;
wire _03297_ ;
wire _03298_ ;
wire _03299_ ;
wire _03300_ ;
wire _03301_ ;
wire _03302_ ;
wire _03303_ ;
wire _03304_ ;
wire _03305_ ;
wire _03306_ ;
wire _03307_ ;
wire _03308_ ;
wire _03309_ ;
wire _03310_ ;
wire _03311_ ;
wire _03312_ ;
wire _03313_ ;
wire _03314_ ;
wire _03315_ ;
wire _03316_ ;
wire _03317_ ;
wire _03318_ ;
wire _03319_ ;
wire _03320_ ;
wire _03321_ ;
wire _03322_ ;
wire _03323_ ;
wire _03324_ ;
wire _03325_ ;
wire _03326_ ;
wire _03327_ ;
wire _03328_ ;
wire _03329_ ;
wire _03330_ ;
wire _03331_ ;
wire _03332_ ;
wire _03333_ ;
wire _03334_ ;
wire _03335_ ;
wire _03336_ ;
wire _03337_ ;
wire _03338_ ;
wire _03339_ ;
wire _03340_ ;
wire _03341_ ;
wire _03342_ ;
wire _03343_ ;
wire _03344_ ;
wire _03345_ ;
wire _03346_ ;
wire _03347_ ;
wire _03348_ ;
wire _03349_ ;
wire _03350_ ;
wire _03351_ ;
wire _03352_ ;
wire _03353_ ;
wire _03354_ ;
wire _03355_ ;
wire _03356_ ;
wire _03357_ ;
wire _03358_ ;
wire _03359_ ;
wire _03360_ ;
wire _03361_ ;
wire _03362_ ;
wire _03363_ ;
wire _03364_ ;
wire _03365_ ;
wire _03366_ ;
wire _03367_ ;
wire _03368_ ;
wire _03369_ ;
wire _03370_ ;
wire _03371_ ;
wire _03372_ ;
wire _03373_ ;
wire _03374_ ;
wire _03375_ ;
wire _03376_ ;
wire _03377_ ;
wire _03378_ ;
wire _03379_ ;
wire _03380_ ;
wire _03381_ ;
wire _03382_ ;
wire _03383_ ;
wire _03384_ ;
wire _03385_ ;
wire _03386_ ;
wire _03387_ ;
wire _03388_ ;
wire _03389_ ;
wire _03390_ ;
wire _03391_ ;
wire _03392_ ;
wire _03393_ ;
wire _03394_ ;
wire _03395_ ;
wire _03396_ ;
wire _03397_ ;
wire _03398_ ;
wire _03399_ ;
wire _03400_ ;
wire _03401_ ;
wire _03402_ ;
wire _03403_ ;
wire _03404_ ;
wire _03405_ ;
wire _03406_ ;
wire _03407_ ;
wire _03408_ ;
wire _03409_ ;
wire _03410_ ;
wire _03411_ ;
wire _03412_ ;
wire _03413_ ;
wire _03414_ ;
wire _03415_ ;
wire _03416_ ;
wire _03417_ ;
wire _03418_ ;
wire _03419_ ;
wire _03420_ ;
wire _03421_ ;
wire _03422_ ;
wire _03423_ ;
wire _03424_ ;
wire _03425_ ;
wire _03426_ ;
wire _03427_ ;
wire _03428_ ;
wire _03429_ ;
wire _03430_ ;
wire _03431_ ;
wire _03432_ ;
wire _03433_ ;
wire _03434_ ;
wire _03435_ ;
wire _03436_ ;
wire _03437_ ;
wire _03438_ ;
wire _03439_ ;
wire _03440_ ;
wire _03441_ ;
wire _03442_ ;
wire _03443_ ;
wire _03444_ ;
wire _03445_ ;
wire _03446_ ;
wire _03447_ ;
wire _03448_ ;
wire _03449_ ;
wire _03450_ ;
wire _03451_ ;
wire _03452_ ;
wire _03453_ ;
wire _03454_ ;
wire _03455_ ;
wire _03456_ ;
wire _03457_ ;
wire _03458_ ;
wire _03459_ ;
wire _03460_ ;
wire _03461_ ;
wire _03462_ ;
wire _03463_ ;
wire _03464_ ;
wire _03465_ ;
wire _03466_ ;
wire _03467_ ;
wire _03468_ ;
wire _03469_ ;
wire _03470_ ;
wire _03471_ ;
wire _03472_ ;
wire _03473_ ;
wire _03474_ ;
wire _03475_ ;
wire _03476_ ;
wire _03477_ ;
wire _03478_ ;
wire _03479_ ;
wire _03480_ ;
wire _03481_ ;
wire _03482_ ;
wire _03483_ ;
wire _03484_ ;
wire _03485_ ;
wire _03486_ ;
wire _03487_ ;
wire _03488_ ;
wire _03489_ ;
wire _03490_ ;
wire _03491_ ;
wire _03492_ ;
wire _03493_ ;
wire _03494_ ;
wire _03495_ ;
wire _03496_ ;
wire _03497_ ;
wire _03498_ ;
wire _03499_ ;
wire _03500_ ;
wire _03501_ ;
wire _03502_ ;
wire _03503_ ;
wire _03504_ ;
wire _03505_ ;
wire _03506_ ;
wire _03507_ ;
wire _03508_ ;
wire _03509_ ;
wire _03510_ ;
wire _03511_ ;
wire _03512_ ;
wire _03513_ ;
wire _03514_ ;
wire _03515_ ;
wire _03516_ ;
wire _03517_ ;
wire _03518_ ;
wire _03519_ ;
wire _03520_ ;
wire _03521_ ;
wire _03522_ ;
wire _03523_ ;
wire _03524_ ;
wire _03525_ ;
wire _03526_ ;
wire _03527_ ;
wire _03528_ ;
wire _03529_ ;
wire _03530_ ;
wire _03531_ ;
wire _03532_ ;
wire _03533_ ;
wire _03534_ ;
wire _03535_ ;
wire _03536_ ;
wire _03537_ ;
wire _03538_ ;
wire _03539_ ;
wire _03540_ ;
wire _03541_ ;
wire _03542_ ;
wire _03543_ ;
wire _03544_ ;
wire _03545_ ;
wire _03546_ ;
wire _03547_ ;
wire _03548_ ;
wire _03549_ ;
wire _03550_ ;
wire _03551_ ;
wire _03552_ ;
wire _03553_ ;
wire _03554_ ;
wire _03555_ ;
wire _03556_ ;
wire _03557_ ;
wire _03558_ ;
wire _03559_ ;
wire _03560_ ;
wire _03561_ ;
wire _03562_ ;
wire _03563_ ;
wire _03564_ ;
wire _03565_ ;
wire _03566_ ;
wire _03567_ ;
wire _03568_ ;
wire _03569_ ;
wire _03570_ ;
wire _03571_ ;
wire _03572_ ;
wire _03573_ ;
wire _03574_ ;
wire _03575_ ;
wire _03576_ ;
wire _03577_ ;
wire _03578_ ;
wire _03579_ ;
wire _03580_ ;
wire _03581_ ;
wire _03582_ ;
wire _03583_ ;
wire _03584_ ;
wire _03585_ ;
wire _03586_ ;
wire _03587_ ;
wire _03588_ ;
wire _03589_ ;
wire _03590_ ;
wire _03591_ ;
wire _03592_ ;
wire _03593_ ;
wire _03594_ ;
wire _03595_ ;
wire _03596_ ;
wire _03597_ ;
wire _03598_ ;
wire _03599_ ;
wire _03600_ ;
wire _03601_ ;
wire _03602_ ;
wire _03603_ ;
wire _03604_ ;
wire _03605_ ;
wire _03606_ ;
wire _03607_ ;
wire _03608_ ;
wire _03609_ ;
wire _03610_ ;
wire _03611_ ;
wire _03612_ ;
wire _03613_ ;
wire _03614_ ;
wire _03615_ ;
wire _03616_ ;
wire _03617_ ;
wire _03618_ ;
wire _03619_ ;
wire _03620_ ;
wire _03621_ ;
wire _03622_ ;
wire _03623_ ;
wire _03624_ ;
wire _03625_ ;
wire _03626_ ;
wire _03627_ ;
wire _03628_ ;
wire _03629_ ;
wire _03630_ ;
wire _03631_ ;
wire _03632_ ;
wire _03633_ ;
wire _03634_ ;
wire _03635_ ;
wire _03636_ ;
wire _03637_ ;
wire _03638_ ;
wire _03639_ ;
wire _03640_ ;
wire _03641_ ;
wire _03642_ ;
wire _03643_ ;
wire _03644_ ;
wire _03645_ ;
wire _03646_ ;
wire _03647_ ;
wire _03648_ ;
wire _03649_ ;
wire _03650_ ;
wire _03651_ ;
wire _03652_ ;
wire _03653_ ;
wire _03654_ ;
wire _03655_ ;
wire _03656_ ;
wire _03657_ ;
wire _03658_ ;
wire _03659_ ;
wire _03660_ ;
wire _03661_ ;
wire _03662_ ;
wire _03663_ ;
wire _03664_ ;
wire _03665_ ;
wire _03666_ ;
wire _03667_ ;
wire _03668_ ;
wire _03669_ ;
wire _03670_ ;
wire _03671_ ;
wire _03672_ ;
wire _03673_ ;
wire _03674_ ;
wire _03675_ ;
wire _03676_ ;
wire _03677_ ;
wire _03678_ ;
wire _03679_ ;
wire _03680_ ;
wire _03681_ ;
wire _03682_ ;
wire _03683_ ;
wire _03684_ ;
wire _03685_ ;
wire _03686_ ;
wire _03687_ ;
wire _03688_ ;
wire _03689_ ;
wire _03690_ ;
wire _03691_ ;
wire _03692_ ;
wire _03693_ ;
wire _03694_ ;
wire _03695_ ;
wire _03696_ ;
wire _03697_ ;
wire _03698_ ;
wire _03699_ ;
wire _03700_ ;
wire _03701_ ;
wire _03702_ ;
wire _03703_ ;
wire _03704_ ;
wire _03705_ ;
wire _03706_ ;
wire _03707_ ;
wire _03708_ ;
wire _03709_ ;
wire _03710_ ;
wire _03711_ ;
wire _03712_ ;
wire _03713_ ;
wire _03714_ ;
wire _03715_ ;
wire _03716_ ;
wire _03717_ ;
wire _03718_ ;
wire _03719_ ;
wire _03720_ ;
wire _03721_ ;
wire _03722_ ;
wire _03723_ ;
wire _03724_ ;
wire _03725_ ;
wire _03726_ ;
wire _03727_ ;
wire _03728_ ;
wire _03729_ ;
wire _03730_ ;
wire _03731_ ;
wire _03732_ ;
wire _03733_ ;
wire _03734_ ;
wire _03735_ ;
wire _03736_ ;
wire _03737_ ;
wire _03738_ ;
wire _03739_ ;
wire _03740_ ;
wire _03741_ ;
wire _03742_ ;
wire _03743_ ;
wire _03744_ ;
wire _03745_ ;
wire _03746_ ;
wire _03747_ ;
wire _03748_ ;
wire _03749_ ;
wire _03750_ ;
wire _03751_ ;
wire _03752_ ;
wire _03753_ ;
wire _03754_ ;
wire _03755_ ;
wire _03756_ ;
wire _03757_ ;
wire _03758_ ;
wire _03759_ ;
wire _03760_ ;
wire _03761_ ;
wire _03762_ ;
wire _03763_ ;
wire _03764_ ;
wire _03765_ ;
wire _03766_ ;
wire _03767_ ;
wire _03768_ ;
wire _03769_ ;
wire _03770_ ;
wire _03771_ ;
wire _03772_ ;
wire _03773_ ;
wire _03774_ ;
wire _03775_ ;
wire _03776_ ;
wire _03777_ ;
wire _03778_ ;
wire _03779_ ;
wire _03780_ ;
wire _03781_ ;
wire _03782_ ;
wire _03783_ ;
wire _03784_ ;
wire _03785_ ;
wire _03786_ ;
wire _03787_ ;
wire _03788_ ;
wire _03789_ ;
wire _03790_ ;
wire _03791_ ;
wire _03792_ ;
wire _03793_ ;
wire _03794_ ;
wire _03795_ ;
wire _03796_ ;
wire _03797_ ;
wire _03798_ ;
wire _03799_ ;
wire _03800_ ;
wire _03801_ ;
wire _03802_ ;
wire _03803_ ;
wire _03804_ ;
wire _03805_ ;
wire _03806_ ;
wire _03807_ ;
wire _03808_ ;
wire _03809_ ;
wire _03810_ ;
wire _03811_ ;
wire _03812_ ;
wire _03813_ ;
wire _03814_ ;
wire _03815_ ;
wire _03816_ ;
wire _03817_ ;
wire _03818_ ;
wire _03819_ ;
wire _03820_ ;
wire _03821_ ;
wire _03822_ ;
wire _03823_ ;
wire _03824_ ;
wire _03825_ ;
wire _03826_ ;
wire _03827_ ;
wire _03828_ ;
wire _03829_ ;
wire _03830_ ;
wire _03831_ ;
wire _03832_ ;
wire _03833_ ;
wire _03834_ ;
wire _03835_ ;
wire _03836_ ;
wire _03837_ ;
wire _03838_ ;
wire _03839_ ;
wire _03840_ ;
wire _03841_ ;
wire _03842_ ;
wire _03843_ ;
wire _03844_ ;
wire _03845_ ;
wire _03846_ ;
wire _03847_ ;
wire _03848_ ;
wire _03849_ ;
wire _03850_ ;
wire _03851_ ;
wire _03852_ ;
wire _03853_ ;
wire _03854_ ;
wire _03855_ ;
wire _03856_ ;
wire _03857_ ;
wire _03858_ ;
wire _03859_ ;
wire _03860_ ;
wire _03861_ ;
wire _03862_ ;
wire _03863_ ;
wire _03864_ ;
wire _03865_ ;
wire _03866_ ;
wire _03867_ ;
wire _03868_ ;
wire _03869_ ;
wire _03870_ ;
wire _03871_ ;
wire _03872_ ;
wire _03873_ ;
wire _03874_ ;
wire _03875_ ;
wire _03876_ ;
wire _03877_ ;
wire _03878_ ;
wire _03879_ ;
wire _03880_ ;
wire _03881_ ;
wire _03882_ ;
wire _03883_ ;
wire _03884_ ;
wire _03885_ ;
wire _03886_ ;
wire _03887_ ;
wire _03888_ ;
wire _03889_ ;
wire _03890_ ;
wire _03891_ ;
wire _03892_ ;
wire _03893_ ;
wire _03894_ ;
wire _03895_ ;
wire _03896_ ;
wire _03897_ ;
wire _03898_ ;
wire _03899_ ;
wire _03900_ ;
wire _03901_ ;
wire _03902_ ;
wire _03903_ ;
wire _03904_ ;
wire _03905_ ;
wire _03906_ ;
wire _03907_ ;
wire _03908_ ;
wire _03909_ ;
wire _03910_ ;
wire _03911_ ;
wire _03912_ ;
wire _03913_ ;
wire _03914_ ;
wire _03915_ ;
wire _03916_ ;
wire _03917_ ;
wire _03918_ ;
wire _03919_ ;
wire _03920_ ;
wire _03921_ ;
wire _03922_ ;
wire _03923_ ;
wire _03924_ ;
wire _03925_ ;
wire _03926_ ;
wire _03927_ ;
wire _03928_ ;
wire _03929_ ;
wire _03930_ ;
wire _03931_ ;
wire _03932_ ;
wire _03933_ ;
wire _03934_ ;
wire _03935_ ;
wire _03936_ ;
wire _03937_ ;
wire _03938_ ;
wire _03939_ ;
wire _03940_ ;
wire _03941_ ;
wire _03942_ ;
wire _03943_ ;
wire _03944_ ;
wire _03945_ ;
wire _03946_ ;
wire _03947_ ;
wire _03948_ ;
wire _03949_ ;
wire _03950_ ;
wire _03951_ ;
wire _03952_ ;
wire _03953_ ;
wire _03954_ ;
wire _03955_ ;
wire _03956_ ;
wire _03957_ ;
wire _03958_ ;
wire _03959_ ;
wire _03960_ ;
wire _03961_ ;
wire _03962_ ;
wire _03963_ ;
wire _03964_ ;
wire _03965_ ;
wire _03966_ ;
wire _03967_ ;
wire _03968_ ;
wire _03969_ ;
wire _03970_ ;
wire _03971_ ;
wire _03972_ ;
wire _03973_ ;
wire _03974_ ;
wire _03975_ ;
wire _03976_ ;
wire _03977_ ;
wire _03978_ ;
wire _03979_ ;
wire _03980_ ;
wire _03981_ ;
wire _03982_ ;
wire _03983_ ;
wire _03984_ ;
wire _03985_ ;
wire _03986_ ;
wire _03987_ ;
wire _03988_ ;
wire _03989_ ;
wire _03990_ ;
wire _03991_ ;
wire _03992_ ;
wire _03993_ ;
wire _03994_ ;
wire _03995_ ;
wire _03996_ ;
wire _03997_ ;
wire _03998_ ;
wire _03999_ ;
wire _04000_ ;
wire _04001_ ;
wire _04002_ ;
wire _04003_ ;
wire _04004_ ;
wire _04005_ ;
wire _04006_ ;
wire _04007_ ;
wire _04008_ ;
wire _04009_ ;
wire _04010_ ;
wire _04011_ ;
wire _04012_ ;
wire _04013_ ;
wire _04014_ ;
wire _04015_ ;
wire _04016_ ;
wire _04017_ ;
wire _04018_ ;
wire _04019_ ;
wire _04020_ ;
wire _04021_ ;
wire _04022_ ;
wire _04023_ ;
wire _04024_ ;
wire _04025_ ;
wire _04026_ ;
wire _04027_ ;
wire _04028_ ;
wire _04029_ ;
wire _04030_ ;
wire _04031_ ;
wire _04032_ ;
wire _04033_ ;
wire _04034_ ;
wire _04035_ ;
wire _04036_ ;
wire _04037_ ;
wire _04038_ ;
wire _04039_ ;
wire _04040_ ;
wire _04041_ ;
wire _04042_ ;
wire _04043_ ;
wire _04044_ ;
wire _04045_ ;
wire _04046_ ;
wire _04047_ ;
wire _04048_ ;
wire _04049_ ;
wire _04050_ ;
wire _04051_ ;
wire _04052_ ;
wire _04053_ ;
wire _04054_ ;
wire _04055_ ;
wire _04056_ ;
wire _04057_ ;
wire _04058_ ;
wire _04059_ ;
wire _04060_ ;
wire _04061_ ;
wire _04062_ ;
wire _04063_ ;
wire _04064_ ;
wire _04065_ ;
wire _04066_ ;
wire _04067_ ;
wire _04068_ ;
wire _04069_ ;
wire _04070_ ;
wire _04071_ ;
wire _04072_ ;
wire _04073_ ;
wire _04074_ ;
wire _04075_ ;
wire _04076_ ;
wire _04077_ ;
wire _04078_ ;
wire _04079_ ;
wire _04080_ ;
wire _04081_ ;
wire _04082_ ;
wire _04083_ ;
wire _04084_ ;
wire _04085_ ;
wire _04086_ ;
wire _04087_ ;
wire _04088_ ;
wire _04089_ ;
wire _04090_ ;
wire _04091_ ;
wire _04092_ ;
wire _04093_ ;
wire _04094_ ;
wire _04095_ ;
wire _04096_ ;
wire _04097_ ;
wire _04098_ ;
wire _04099_ ;
wire _04100_ ;
wire _04101_ ;
wire _04102_ ;
wire _04103_ ;
wire _04104_ ;
wire _04105_ ;
wire _04106_ ;
wire _04107_ ;
wire _04108_ ;
wire _04109_ ;
wire _04110_ ;
wire _04111_ ;
wire _04112_ ;
wire _04113_ ;
wire _04114_ ;
wire _04115_ ;
wire _04116_ ;
wire _04117_ ;
wire _04118_ ;
wire _04119_ ;
wire _04120_ ;
wire _04121_ ;
wire _04122_ ;
wire _04123_ ;
wire _04124_ ;
wire _04125_ ;
wire _04126_ ;
wire _04127_ ;
wire _04128_ ;
wire _04129_ ;
wire _04130_ ;
wire _04131_ ;
wire _04132_ ;
wire _04133_ ;
wire _04134_ ;
wire _04135_ ;
wire _04136_ ;
wire _04137_ ;
wire _04138_ ;
wire _04139_ ;
wire _04140_ ;
wire _04141_ ;
wire _04142_ ;
wire _04143_ ;
wire _04144_ ;
wire _04145_ ;
wire _04146_ ;
wire _04147_ ;
wire _04148_ ;
wire _04149_ ;
wire _04150_ ;
wire _04151_ ;
wire _04152_ ;
wire _04153_ ;
wire _04154_ ;
wire _04155_ ;
wire _04156_ ;
wire _04157_ ;
wire _04158_ ;
wire _04159_ ;
wire _04160_ ;
wire _04161_ ;
wire _04162_ ;
wire _04163_ ;
wire _04164_ ;
wire _04165_ ;
wire _04166_ ;
wire _04167_ ;
wire _04168_ ;
wire _04169_ ;
wire _04170_ ;
wire _04171_ ;
wire _04172_ ;
wire _04173_ ;
wire _04174_ ;
wire _04175_ ;
wire _04176_ ;
wire _04177_ ;
wire _04178_ ;
wire _04179_ ;
wire _04180_ ;
wire _04181_ ;
wire _04182_ ;
wire _04183_ ;
wire _04184_ ;
wire _04185_ ;
wire _04186_ ;
wire _04187_ ;
wire _04188_ ;
wire _04189_ ;
wire _04190_ ;
wire _04191_ ;
wire _04192_ ;
wire _04193_ ;
wire _04194_ ;
wire _04195_ ;
wire _04196_ ;
wire _04197_ ;
wire _04198_ ;
wire _04199_ ;
wire _04200_ ;
wire _04201_ ;
wire _04202_ ;
wire _04203_ ;
wire _04204_ ;
wire _04205_ ;
wire _04206_ ;
wire _04207_ ;
wire _04208_ ;
wire _04209_ ;
wire _04210_ ;
wire _04211_ ;
wire _04212_ ;
wire _04213_ ;
wire _04214_ ;
wire _04215_ ;
wire _04216_ ;
wire _04217_ ;
wire _04218_ ;
wire _04219_ ;
wire _04220_ ;
wire _04221_ ;
wire _04222_ ;
wire _04223_ ;
wire _04224_ ;
wire _04225_ ;
wire _04226_ ;
wire _04227_ ;
wire _04228_ ;
wire _04229_ ;
wire _04230_ ;
wire _04231_ ;
wire _04232_ ;
wire _04233_ ;
wire _04234_ ;
wire _04235_ ;
wire _04236_ ;
wire _04237_ ;
wire _04238_ ;
wire _04239_ ;
wire _04240_ ;
wire _04241_ ;
wire _04242_ ;
wire _04243_ ;
wire _04244_ ;
wire _04245_ ;
wire _04246_ ;
wire _04247_ ;
wire _04248_ ;
wire _04249_ ;
wire _04250_ ;
wire _04251_ ;
wire _04252_ ;
wire _04253_ ;
wire _04254_ ;
wire _04255_ ;
wire _04256_ ;
wire _04257_ ;
wire _04258_ ;
wire _04259_ ;
wire _04260_ ;
wire _04261_ ;
wire _04262_ ;
wire _04263_ ;
wire _04264_ ;
wire _04265_ ;
wire _04266_ ;
wire _04267_ ;
wire _04268_ ;
wire _04269_ ;
wire _04270_ ;
wire _04271_ ;
wire _04272_ ;
wire _04273_ ;
wire _04274_ ;
wire _04275_ ;
wire _04276_ ;
wire _04277_ ;
wire _04278_ ;
wire _04279_ ;
wire _04280_ ;
wire _04281_ ;
wire _04282_ ;
wire _04283_ ;
wire _04284_ ;
wire _04285_ ;
wire _04286_ ;
wire _04287_ ;
wire _04288_ ;
wire _04289_ ;
wire _04290_ ;
wire _04291_ ;
wire _04292_ ;
wire _04293_ ;
wire _04294_ ;
wire _04295_ ;
wire _04296_ ;
wire _04297_ ;
wire _04298_ ;
wire _04299_ ;
wire _04300_ ;
wire _04301_ ;
wire _04302_ ;
wire _04303_ ;
wire _04304_ ;
wire _04305_ ;
wire _04306_ ;
wire _04307_ ;
wire _04308_ ;
wire _04309_ ;
wire _04310_ ;
wire _04311_ ;
wire _04312_ ;
wire _04313_ ;
wire _04314_ ;
wire _04315_ ;
wire _04316_ ;
wire _04317_ ;
wire _04318_ ;
wire _04319_ ;
wire _04320_ ;
wire _04321_ ;
wire _04322_ ;
wire _04323_ ;
wire _04324_ ;
wire _04325_ ;
wire _04326_ ;
wire _04327_ ;
wire _04328_ ;
wire _04329_ ;
wire _04330_ ;
wire _04331_ ;
wire _04332_ ;
wire _04333_ ;
wire _04334_ ;
wire _04335_ ;
wire _04336_ ;
wire _04337_ ;
wire _04338_ ;
wire _04339_ ;
wire _04340_ ;
wire _04341_ ;
wire _04342_ ;
wire _04343_ ;
wire _04344_ ;
wire _04345_ ;
wire _04346_ ;
wire _04347_ ;
wire _04348_ ;
wire _04349_ ;
wire _04350_ ;
wire _04351_ ;
wire _04352_ ;
wire _04353_ ;
wire _04354_ ;
wire _04355_ ;
wire _04356_ ;
wire _04357_ ;
wire _04358_ ;
wire _04359_ ;
wire _04360_ ;
wire _04361_ ;
wire _04362_ ;
wire _04363_ ;
wire _04364_ ;
wire _04365_ ;
wire _04366_ ;
wire _04367_ ;
wire _04368_ ;
wire _04369_ ;
wire _04370_ ;
wire _04371_ ;
wire _04372_ ;
wire _04373_ ;
wire _04374_ ;
wire _04375_ ;
wire _04376_ ;
wire _04377_ ;
wire _04378_ ;
wire _04379_ ;
wire _04380_ ;
wire _04381_ ;
wire _04382_ ;
wire _04383_ ;
wire _04384_ ;
wire _04385_ ;
wire _04386_ ;
wire _04387_ ;
wire _04388_ ;
wire _04389_ ;
wire _04390_ ;
wire _04391_ ;
wire _04392_ ;
wire _04393_ ;
wire _04394_ ;
wire _04395_ ;
wire _04396_ ;
wire _04397_ ;
wire _04398_ ;
wire _04399_ ;
wire _04400_ ;
wire _04401_ ;
wire _04402_ ;
wire _04403_ ;
wire _04404_ ;
wire _04405_ ;
wire _04406_ ;
wire _04407_ ;
wire _04408_ ;
wire _04409_ ;
wire _04410_ ;
wire _04411_ ;
wire _04412_ ;
wire _04413_ ;
wire _04414_ ;
wire _04415_ ;
wire _04416_ ;
wire _04417_ ;
wire _04418_ ;
wire _04419_ ;
wire _04420_ ;
wire _04421_ ;
wire _04422_ ;
wire _04423_ ;
wire _04424_ ;
wire _04425_ ;
wire _04426_ ;
wire _04427_ ;
wire _04428_ ;
wire _04429_ ;
wire _04430_ ;
wire _04431_ ;
wire _04432_ ;
wire _04433_ ;
wire _04434_ ;
wire _04435_ ;
wire _04436_ ;
wire _04437_ ;
wire _04438_ ;
wire _04439_ ;
wire _04440_ ;
wire _04441_ ;
wire _04442_ ;
wire _04443_ ;
wire _04444_ ;
wire _04445_ ;
wire _04446_ ;
wire _04447_ ;
wire _04448_ ;
wire _04449_ ;
wire _04450_ ;
wire _04451_ ;
wire _04452_ ;
wire _04453_ ;
wire _04454_ ;
wire _04455_ ;
wire _04456_ ;
wire _04457_ ;
wire _04458_ ;
wire _04459_ ;
wire _04460_ ;
wire _04461_ ;
wire _04462_ ;
wire _04463_ ;
wire _04464_ ;
wire _04465_ ;
wire _04466_ ;
wire _04467_ ;
wire _04468_ ;
wire _04469_ ;
wire _04470_ ;
wire _04471_ ;
wire _04472_ ;
wire _04473_ ;
wire _04474_ ;
wire _04475_ ;
wire _04476_ ;
wire _04477_ ;
wire _04478_ ;
wire _04479_ ;
wire _04480_ ;
wire _04481_ ;
wire _04482_ ;
wire _04483_ ;
wire _04484_ ;
wire _04485_ ;
wire _04486_ ;
wire _04487_ ;
wire _04488_ ;
wire _04489_ ;
wire _04490_ ;
wire _04491_ ;
wire _04492_ ;
wire _04493_ ;
wire _04494_ ;
wire _04495_ ;
wire _04496_ ;
wire _04497_ ;
wire _04498_ ;
wire _04499_ ;
wire _04500_ ;
wire _04501_ ;
wire _04502_ ;
wire _04503_ ;
wire _04504_ ;
wire _04505_ ;
wire _04506_ ;
wire _04507_ ;
wire _04508_ ;
wire _04509_ ;
wire _04510_ ;
wire _04511_ ;
wire _04512_ ;
wire _04513_ ;
wire _04514_ ;
wire _04515_ ;
wire _04516_ ;
wire _04517_ ;
wire _04518_ ;
wire _04519_ ;
wire _04520_ ;
wire _04521_ ;
wire _04522_ ;
wire _04523_ ;
wire _04524_ ;
wire _04525_ ;
wire _04526_ ;
wire _04527_ ;
wire _04528_ ;
wire _04529_ ;
wire _04530_ ;
wire _04531_ ;
wire _04532_ ;
wire _04533_ ;
wire _04534_ ;
wire _04535_ ;
wire _04536_ ;
wire _04537_ ;
wire _04538_ ;
wire _04539_ ;
wire _04540_ ;
wire _04541_ ;
wire _04542_ ;
wire _04543_ ;
wire _04544_ ;
wire _04545_ ;
wire _04546_ ;
wire _04547_ ;
wire _04548_ ;
wire _04549_ ;
wire _04550_ ;
wire _04551_ ;
wire _04552_ ;
wire _04553_ ;
wire _04554_ ;
wire _04555_ ;
wire _04556_ ;
wire _04557_ ;
wire _04558_ ;
wire _04559_ ;
wire _04560_ ;
wire _04561_ ;
wire _04562_ ;
wire _04563_ ;
wire _04564_ ;
wire _04565_ ;
wire _04566_ ;
wire _04567_ ;
wire _04568_ ;
wire _04569_ ;
wire _04570_ ;
wire _04571_ ;
wire _04572_ ;
wire _04573_ ;
wire _04574_ ;
wire _04575_ ;
wire _04576_ ;
wire _04577_ ;
wire _04578_ ;
wire _04579_ ;
wire _04580_ ;
wire _04581_ ;
wire _04582_ ;
wire _04583_ ;
wire _04584_ ;
wire _04585_ ;
wire _04586_ ;
wire _04587_ ;
wire _04588_ ;
wire _04589_ ;
wire _04590_ ;
wire _04591_ ;
wire _04592_ ;
wire _04593_ ;
wire _04594_ ;
wire _04595_ ;
wire _04596_ ;
wire _04597_ ;
wire _04598_ ;
wire _04599_ ;
wire _04600_ ;
wire _04601_ ;
wire _04602_ ;
wire _04603_ ;
wire _04604_ ;
wire _04605_ ;
wire _04606_ ;
wire _04607_ ;
wire _04608_ ;
wire _04609_ ;
wire _04610_ ;
wire _04611_ ;
wire _04612_ ;
wire _04613_ ;
wire _04614_ ;
wire _04615_ ;
wire _04616_ ;
wire _04617_ ;
wire _04618_ ;
wire _04619_ ;
wire _04620_ ;
wire _04621_ ;
wire _04622_ ;
wire _04623_ ;
wire _04624_ ;
wire _04625_ ;
wire _04626_ ;
wire _04627_ ;
wire _04628_ ;
wire _04629_ ;
wire _04630_ ;
wire _04631_ ;
wire _04632_ ;
wire _04633_ ;
wire _04634_ ;
wire _04635_ ;
wire _04636_ ;
wire _04637_ ;
wire _04638_ ;
wire _04639_ ;
wire _04640_ ;
wire _04641_ ;
wire _04642_ ;
wire _04643_ ;
wire _04644_ ;
wire _04645_ ;
wire _04646_ ;
wire _04647_ ;
wire _04648_ ;
wire _04649_ ;
wire _04650_ ;
wire _04651_ ;
wire _04652_ ;
wire _04653_ ;
wire _04654_ ;
wire _04655_ ;
wire _04656_ ;
wire _04657_ ;
wire _04658_ ;
wire _04659_ ;
wire _04660_ ;
wire _04661_ ;
wire _04662_ ;
wire _04663_ ;
wire _04664_ ;
wire _04665_ ;
wire _04666_ ;
wire _04667_ ;
wire _04668_ ;
wire _04669_ ;
wire _04670_ ;
wire _04671_ ;
wire _04672_ ;
wire _04673_ ;
wire _04674_ ;
wire _04675_ ;
wire _04676_ ;
wire _04677_ ;
wire _04678_ ;
wire _04679_ ;
wire _04680_ ;
wire _04681_ ;
wire _04682_ ;
wire _04683_ ;
wire _04684_ ;
wire _04685_ ;
wire _04686_ ;
wire _04687_ ;
wire _04688_ ;
wire _04689_ ;
wire _04690_ ;
wire _04691_ ;
wire _04692_ ;
wire _04693_ ;
wire _04694_ ;
wire _04695_ ;
wire _04696_ ;
wire _04697_ ;
wire _04698_ ;
wire _04699_ ;
wire _04700_ ;
wire _04701_ ;
wire _04702_ ;
wire _04703_ ;
wire _04704_ ;
wire _04705_ ;
wire _04706_ ;
wire _04707_ ;
wire _04708_ ;
wire _04709_ ;
wire _04710_ ;
wire _04711_ ;
wire _04712_ ;
wire _04713_ ;
wire _04714_ ;
wire _04715_ ;
wire _04716_ ;
wire _04717_ ;
wire _04718_ ;
wire _04719_ ;
wire _04720_ ;
wire _04721_ ;
wire _04722_ ;
wire _04723_ ;
wire _04724_ ;
wire _04725_ ;
wire _04726_ ;
wire _04727_ ;
wire _04728_ ;
wire _04729_ ;
wire _04730_ ;
wire _04731_ ;
wire _04732_ ;
wire _04733_ ;
wire _04734_ ;
wire _04735_ ;
wire _04736_ ;
wire _04737_ ;
wire _04738_ ;
wire _04739_ ;
wire _04740_ ;
wire _04741_ ;
wire _04742_ ;
wire _04743_ ;
wire _04744_ ;
wire _04745_ ;
wire _04746_ ;
wire _04747_ ;
wire _04748_ ;
wire _04749_ ;
wire _04750_ ;
wire _04751_ ;
wire _04752_ ;
wire _04753_ ;
wire _04754_ ;
wire _04755_ ;
wire _04756_ ;
wire _04757_ ;
wire _04758_ ;
wire _04759_ ;
wire _04760_ ;
wire _04761_ ;
wire _04762_ ;
wire _04763_ ;
wire _04764_ ;
wire _04765_ ;
wire _04766_ ;
wire _04767_ ;
wire _04768_ ;
wire _04769_ ;
wire _04770_ ;
wire _04771_ ;
wire _04772_ ;
wire _04773_ ;
wire _04774_ ;
wire _04775_ ;
wire _04776_ ;
wire _04777_ ;
wire _04778_ ;
wire _04779_ ;
wire _04780_ ;
wire _04781_ ;
wire _04782_ ;
wire _04783_ ;
wire _04784_ ;
wire _04785_ ;
wire _04786_ ;
wire _04787_ ;
wire _04788_ ;
wire _04789_ ;
wire _04790_ ;
wire _04791_ ;
wire _04792_ ;
wire _04793_ ;
wire _04794_ ;
wire _04795_ ;
wire _04796_ ;
wire _04797_ ;
wire _04798_ ;
wire _04799_ ;
wire _04800_ ;
wire _04801_ ;
wire _04802_ ;
wire _04803_ ;
wire _04804_ ;
wire _04805_ ;
wire _04806_ ;
wire _04807_ ;
wire _04808_ ;
wire _04809_ ;
wire _04810_ ;
wire _04811_ ;
wire _04812_ ;
wire _04813_ ;
wire _04814_ ;
wire _04815_ ;
wire _04816_ ;
wire _04817_ ;
wire _04818_ ;
wire _04819_ ;
wire _04820_ ;
wire _04821_ ;
wire _04822_ ;
wire _04823_ ;
wire _04824_ ;
wire _04825_ ;
wire _04826_ ;
wire _04827_ ;
wire _04828_ ;
wire _04829_ ;
wire _04830_ ;
wire _04831_ ;
wire _04832_ ;
wire _04833_ ;
wire _04834_ ;
wire _04835_ ;
wire _04836_ ;
wire _04837_ ;
wire _04838_ ;
wire _04839_ ;
wire _04840_ ;
wire _04841_ ;
wire _04842_ ;
wire _04843_ ;
wire _04844_ ;
wire _04845_ ;
wire _04846_ ;
wire _04847_ ;
wire _04848_ ;
wire _04849_ ;
wire _04850_ ;
wire _04851_ ;
wire _04852_ ;
wire _04853_ ;
wire _04854_ ;
wire _04855_ ;
wire _04856_ ;
wire _04857_ ;
wire _04858_ ;
wire _04859_ ;
wire _04860_ ;
wire _04861_ ;
wire _04862_ ;
wire _04863_ ;
wire _04864_ ;
wire _04865_ ;
wire _04866_ ;
wire _04867_ ;
wire _04868_ ;
wire _04869_ ;
wire _04870_ ;
wire _04871_ ;
wire _04872_ ;
wire _04873_ ;
wire _04874_ ;
wire _04875_ ;
wire _04876_ ;
wire _04877_ ;
wire _04878_ ;
wire _04879_ ;
wire _04880_ ;
wire _04881_ ;
wire _04882_ ;
wire _04883_ ;
wire _04884_ ;
wire _04885_ ;
wire _04886_ ;
wire _04887_ ;
wire _04888_ ;
wire _04889_ ;
wire _04890_ ;
wire _04891_ ;
wire _04892_ ;
wire _04893_ ;
wire _04894_ ;
wire _04895_ ;
wire _04896_ ;
wire _04897_ ;
wire _04898_ ;
wire _04899_ ;
wire _04900_ ;
wire _04901_ ;
wire _04902_ ;
wire _04903_ ;
wire _04904_ ;
wire _04905_ ;
wire _04906_ ;
wire _04907_ ;
wire _04908_ ;
wire _04909_ ;
wire _04910_ ;
wire _04911_ ;
wire _04912_ ;
wire _04913_ ;
wire _04914_ ;
wire _04915_ ;
wire _04916_ ;
wire _04917_ ;
wire _04918_ ;
wire _04919_ ;
wire _04920_ ;
wire _04921_ ;
wire _04922_ ;
wire _04923_ ;
wire _04924_ ;
wire _04925_ ;
wire _04926_ ;
wire _04927_ ;
wire _04928_ ;
wire _04929_ ;
wire _04930_ ;
wire _04931_ ;
wire _04932_ ;
wire _04933_ ;
wire _04934_ ;
wire _04935_ ;
wire _04936_ ;
wire _04937_ ;
wire _04938_ ;
wire _04939_ ;
wire _04940_ ;
wire _04941_ ;
wire _04942_ ;
wire _04943_ ;
wire _04944_ ;
wire _04945_ ;
wire _04946_ ;
wire _04947_ ;
wire _04948_ ;
wire _04949_ ;
wire _04950_ ;
wire _04951_ ;
wire _04952_ ;
wire _04953_ ;
wire _04954_ ;
wire _04955_ ;
wire _04956_ ;
wire _04957_ ;
wire _04958_ ;
wire _04959_ ;
wire _04960_ ;
wire _04961_ ;
wire _04962_ ;
wire _04963_ ;
wire _04964_ ;
wire _04965_ ;
wire _04966_ ;
wire _04967_ ;
wire _04968_ ;
wire _04969_ ;
wire _04970_ ;
wire _04971_ ;
wire _04972_ ;
wire _04973_ ;
wire _04974_ ;
wire _04975_ ;
wire _04976_ ;
wire _04977_ ;
wire _04978_ ;
wire _04979_ ;
wire _04980_ ;
wire _04981_ ;
wire _04982_ ;
wire _04983_ ;
wire _04984_ ;
wire _04985_ ;
wire _04986_ ;
wire _04987_ ;
wire _04988_ ;
wire _04989_ ;
wire _04990_ ;
wire _04991_ ;
wire _04992_ ;
wire _04993_ ;
wire _04994_ ;
wire _04995_ ;
wire _04996_ ;
wire _04997_ ;
wire _04998_ ;
wire _04999_ ;
wire _05000_ ;
wire _05001_ ;
wire _05002_ ;
wire _05003_ ;
wire _05004_ ;
wire _05005_ ;
wire _05006_ ;
wire _05007_ ;
wire _05008_ ;
wire _05009_ ;
wire _05010_ ;
wire _05011_ ;
wire _05012_ ;
wire _05013_ ;
wire _05014_ ;
wire _05015_ ;
wire _05016_ ;
wire _05017_ ;
wire _05018_ ;
wire _05019_ ;
wire _05020_ ;
wire _05021_ ;
wire _05022_ ;
wire _05023_ ;
wire _05024_ ;
wire _05025_ ;
wire _05026_ ;
wire _05027_ ;
wire _05028_ ;
wire _05029_ ;
wire _05030_ ;
wire _05031_ ;
wire _05032_ ;
wire _05033_ ;
wire _05034_ ;
wire _05035_ ;
wire _05036_ ;
wire _05037_ ;
wire _05038_ ;
wire _05039_ ;
wire _05040_ ;
wire _05041_ ;
wire _05042_ ;
wire _05043_ ;
wire _05044_ ;
wire _05045_ ;
wire _05046_ ;
wire _05047_ ;
wire _05048_ ;
wire _05049_ ;
wire _05050_ ;
wire _05051_ ;
wire _05052_ ;
wire _05053_ ;
wire _05054_ ;
wire _05055_ ;
wire _05056_ ;
wire _05057_ ;
wire _05058_ ;
wire _05059_ ;
wire _05060_ ;
wire _05061_ ;
wire _05062_ ;
wire _05063_ ;
wire _05064_ ;
wire _05065_ ;
wire _05066_ ;
wire _05067_ ;
wire _05068_ ;
wire _05069_ ;
wire _05070_ ;
wire _05071_ ;
wire _05072_ ;
wire _05073_ ;
wire _05074_ ;
wire _05075_ ;
wire _05076_ ;
wire _05077_ ;
wire _05078_ ;
wire _05079_ ;
wire _05080_ ;
wire _05081_ ;
wire _05082_ ;
wire _05083_ ;
wire _05084_ ;
wire _05085_ ;
wire _05086_ ;
wire _05087_ ;
wire _05088_ ;
wire _05089_ ;
wire _05090_ ;
wire _05091_ ;
wire _05092_ ;
wire _05093_ ;
wire _05094_ ;
wire _05095_ ;
wire _05096_ ;
wire _05097_ ;
wire _05098_ ;
wire _05099_ ;
wire _05100_ ;
wire _05101_ ;
wire _05102_ ;
wire _05103_ ;
wire _05104_ ;
wire _05105_ ;
wire _05106_ ;
wire _05107_ ;
wire _05108_ ;
wire _05109_ ;
wire _05110_ ;
wire _05111_ ;
wire _05112_ ;
wire _05113_ ;
wire _05114_ ;
wire _05115_ ;
wire _05116_ ;
wire _05117_ ;
wire _05118_ ;
wire _05119_ ;
wire _05120_ ;
wire _05121_ ;
wire _05122_ ;
wire _05123_ ;
wire _05124_ ;
wire _05125_ ;
wire _05126_ ;
wire _05127_ ;
wire _05128_ ;
wire _05129_ ;
wire _05130_ ;
wire _05131_ ;
wire _05132_ ;
wire _05133_ ;
wire _05134_ ;
wire _05135_ ;
wire _05136_ ;
wire _05137_ ;
wire _05138_ ;
wire _05139_ ;
wire _05140_ ;
wire _05141_ ;
wire _05142_ ;
wire _05143_ ;
wire _05144_ ;
wire _05145_ ;
wire _05146_ ;
wire _05147_ ;
wire _05148_ ;
wire _05149_ ;
wire _05150_ ;
wire _05151_ ;
wire _05152_ ;
wire _05153_ ;
wire _05154_ ;
wire _05155_ ;
wire _05156_ ;
wire _05157_ ;
wire _05158_ ;
wire _05159_ ;
wire _05160_ ;
wire _05161_ ;
wire _05162_ ;
wire _05163_ ;
wire _05164_ ;
wire _05165_ ;
wire _05166_ ;
wire _05167_ ;
wire _05168_ ;
wire _05169_ ;
wire _05170_ ;
wire _05171_ ;
wire _05172_ ;
wire _05173_ ;
wire _05174_ ;
wire _05175_ ;
wire _05176_ ;
wire _05177_ ;
wire _05178_ ;
wire _05179_ ;
wire _05180_ ;
wire _05181_ ;
wire _05182_ ;
wire _05183_ ;
wire _05184_ ;
wire _05185_ ;
wire _05186_ ;
wire _05187_ ;
wire _05188_ ;
wire _05189_ ;
wire _05190_ ;
wire _05191_ ;
wire _05192_ ;
wire _05193_ ;
wire _05194_ ;
wire _05195_ ;
wire _05196_ ;
wire _05197_ ;
wire _05198_ ;
wire _05199_ ;
wire _05200_ ;
wire _05201_ ;
wire _05202_ ;
wire _05203_ ;
wire _05204_ ;
wire _05205_ ;
wire _05206_ ;
wire _05207_ ;
wire _05208_ ;
wire _05209_ ;
wire _05210_ ;
wire _05211_ ;
wire _05212_ ;
wire _05213_ ;
wire _05214_ ;
wire _05215_ ;
wire _05216_ ;
wire _05217_ ;
wire _05218_ ;
wire _05219_ ;
wire _05220_ ;
wire _05221_ ;
wire _05222_ ;
wire _05223_ ;
wire _05224_ ;
wire _05225_ ;
wire _05226_ ;
wire _05227_ ;
wire _05228_ ;
wire _05229_ ;
wire _05230_ ;
wire _05231_ ;
wire _05232_ ;
wire _05233_ ;
wire _05234_ ;
wire _05235_ ;
wire _05236_ ;
wire _05237_ ;
wire _05238_ ;
wire _05239_ ;
wire _05240_ ;
wire _05241_ ;
wire _05242_ ;
wire _05243_ ;
wire _05244_ ;
wire _05245_ ;
wire _05246_ ;
wire _05247_ ;
wire _05248_ ;
wire _05249_ ;
wire _05250_ ;
wire _05251_ ;
wire _05252_ ;
wire _05253_ ;
wire _05254_ ;
wire _05255_ ;
wire _05256_ ;
wire _05257_ ;
wire _05258_ ;
wire _05259_ ;
wire _05260_ ;
wire _05261_ ;
wire _05262_ ;
wire _05263_ ;
wire _05264_ ;
wire _05265_ ;
wire _05266_ ;
wire _05267_ ;
wire _05268_ ;
wire _05269_ ;
wire _05270_ ;
wire _05271_ ;
wire _05272_ ;
wire _05273_ ;
wire _05274_ ;
wire _05275_ ;
wire _05276_ ;
wire _05277_ ;
wire _05278_ ;
wire _05279_ ;
wire _05280_ ;
wire _05281_ ;
wire _05282_ ;
wire _05283_ ;
wire _05284_ ;
wire _05285_ ;
wire _05286_ ;
wire _05287_ ;
wire _05288_ ;
wire _05289_ ;
wire _05290_ ;
wire _05291_ ;
wire _05292_ ;
wire _05293_ ;
wire _05294_ ;
wire _05295_ ;
wire _05296_ ;
wire _05297_ ;
wire _05298_ ;
wire _05299_ ;
wire _05300_ ;
wire _05301_ ;
wire _05302_ ;
wire _05303_ ;
wire _05304_ ;
wire _05305_ ;
wire _05306_ ;
wire _05307_ ;
wire _05308_ ;
wire _05309_ ;
wire _05310_ ;
wire _05311_ ;
wire _05312_ ;
wire _05313_ ;
wire _05314_ ;
wire _05315_ ;
wire _05316_ ;
wire _05317_ ;
wire _05318_ ;
wire _05319_ ;
wire _05320_ ;
wire _05321_ ;
wire _05322_ ;
wire _05323_ ;
wire _05324_ ;
wire _05325_ ;
wire _05326_ ;
wire _05327_ ;
wire _05328_ ;
wire _05329_ ;
wire _05330_ ;
wire _05331_ ;
wire _05332_ ;
wire _05333_ ;
wire _05334_ ;
wire _05335_ ;
wire _05336_ ;
wire _05337_ ;
wire _05338_ ;
wire _05339_ ;
wire _05340_ ;
wire _05341_ ;
wire _05342_ ;
wire _05343_ ;
wire _05344_ ;
wire _05345_ ;
wire _05346_ ;
wire _05347_ ;
wire _05348_ ;
wire _05349_ ;
wire _05350_ ;
wire _05351_ ;
wire _05352_ ;
wire _05353_ ;
wire _05354_ ;
wire _05355_ ;
wire _05356_ ;
wire _05357_ ;
wire _05358_ ;
wire _05359_ ;
wire _05360_ ;
wire _05361_ ;
wire _05362_ ;
wire _05363_ ;
wire _05364_ ;
wire _05365_ ;
wire _05366_ ;
wire _05367_ ;
wire _05368_ ;
wire _05369_ ;
wire _05370_ ;
wire _05371_ ;
wire _05372_ ;
wire _05373_ ;
wire _05374_ ;
wire _05375_ ;
wire _05376_ ;
wire _05377_ ;
wire _05378_ ;
wire _05379_ ;
wire _05380_ ;
wire _05381_ ;
wire _05382_ ;
wire _05383_ ;
wire _05384_ ;
wire _05385_ ;
wire _05386_ ;
wire _05387_ ;
wire _05388_ ;
wire _05389_ ;
wire _05390_ ;
wire _05391_ ;
wire _05392_ ;
wire _05393_ ;
wire _05394_ ;
wire _05395_ ;
wire _05396_ ;
wire _05397_ ;
wire _05398_ ;
wire _05399_ ;
wire _05400_ ;
wire _05401_ ;
wire _05402_ ;
wire _05403_ ;
wire _05404_ ;
wire _05405_ ;
wire _05406_ ;
wire _05407_ ;
wire _05408_ ;
wire _05409_ ;
wire _05410_ ;
wire _05411_ ;
wire _05412_ ;
wire _05413_ ;
wire _05414_ ;
wire _05415_ ;
wire _05416_ ;
wire _05417_ ;
wire _05418_ ;
wire _05419_ ;
wire _05420_ ;
wire _05421_ ;
wire _05422_ ;
wire _05423_ ;
wire _05424_ ;
wire _05425_ ;
wire _05426_ ;
wire _05427_ ;
wire _05428_ ;
wire _05429_ ;
wire _05430_ ;
wire _05431_ ;
wire _05432_ ;
wire _05433_ ;
wire _05434_ ;
wire _05435_ ;
wire _05436_ ;
wire _05437_ ;
wire _05438_ ;
wire _05439_ ;
wire _05440_ ;
wire _05441_ ;
wire _05442_ ;
wire _05443_ ;
wire _05444_ ;
wire _05445_ ;
wire _05446_ ;
wire _05447_ ;
wire _05448_ ;
wire _05449_ ;
wire _05450_ ;
wire _05451_ ;
wire _05452_ ;
wire _05453_ ;
wire _05454_ ;
wire _05455_ ;
wire _05456_ ;
wire _05457_ ;
wire _05458_ ;
wire _05459_ ;
wire _05460_ ;
wire _05461_ ;
wire _05462_ ;
wire _05463_ ;
wire _05464_ ;
wire _05465_ ;
wire _05466_ ;
wire _05467_ ;
wire _05468_ ;
wire _05469_ ;
wire _05470_ ;
wire _05471_ ;
wire _05472_ ;
wire _05473_ ;
wire _05474_ ;
wire _05475_ ;
wire _05476_ ;
wire _05477_ ;
wire _05478_ ;
wire _05479_ ;
wire _05480_ ;
wire _05481_ ;
wire _05482_ ;
wire _05483_ ;
wire _05484_ ;
wire _05485_ ;
wire _05486_ ;
wire _05487_ ;
wire _05488_ ;
wire _05489_ ;
wire _05490_ ;
wire _05491_ ;
wire _05492_ ;
wire _05493_ ;
wire _05494_ ;
wire _05495_ ;
wire _05496_ ;
wire _05497_ ;
wire _05498_ ;
wire _05499_ ;
wire _05500_ ;
wire _05501_ ;
wire _05502_ ;
wire _05503_ ;
wire _05504_ ;
wire _05505_ ;
wire _05506_ ;
wire _05507_ ;
wire _05508_ ;
wire _05509_ ;
wire _05510_ ;
wire _05511_ ;
wire _05512_ ;
wire _05513_ ;
wire _05514_ ;
wire _05515_ ;
wire _05516_ ;
wire _05517_ ;
wire _05518_ ;
wire _05519_ ;
wire _05520_ ;
wire _05521_ ;
wire _05522_ ;
wire _05523_ ;
wire _05524_ ;
wire _05525_ ;
wire _05526_ ;
wire _05527_ ;
wire _05528_ ;
wire _05529_ ;
wire _05530_ ;
wire _05531_ ;
wire _05532_ ;
wire _05533_ ;
wire _05534_ ;
wire _05535_ ;
wire _05536_ ;
wire _05537_ ;
wire _05538_ ;
wire _05539_ ;
wire _05540_ ;
wire _05541_ ;
wire _05542_ ;
wire _05543_ ;
wire _05544_ ;
wire _05545_ ;
wire _05546_ ;
wire _05547_ ;
wire _05548_ ;
wire _05549_ ;
wire _05550_ ;
wire _05551_ ;
wire _05552_ ;
wire _05553_ ;
wire _05554_ ;
wire _05555_ ;
wire _05556_ ;
wire _05557_ ;
wire _05558_ ;
wire _05559_ ;
wire _05560_ ;
wire _05561_ ;
wire _05562_ ;
wire _05563_ ;
wire _05564_ ;
wire _05565_ ;
wire _05566_ ;
wire _05567_ ;
wire _05568_ ;
wire _05569_ ;
wire _05570_ ;
wire _05571_ ;
wire _05572_ ;
wire _05573_ ;
wire _05574_ ;
wire _05575_ ;
wire _05576_ ;
wire _05577_ ;
wire _05578_ ;
wire _05579_ ;
wire _05580_ ;
wire _05581_ ;
wire _05582_ ;
wire _05583_ ;
wire _05584_ ;
wire _05585_ ;
wire _05586_ ;
wire _05587_ ;
wire _05588_ ;
wire _05589_ ;
wire _05590_ ;
wire _05591_ ;
wire _05592_ ;
wire _05593_ ;
wire _05594_ ;
wire _05595_ ;
wire _05596_ ;
wire _05597_ ;
wire _05598_ ;
wire _05599_ ;
wire _05600_ ;
wire _05601_ ;
wire _05602_ ;
wire _05603_ ;
wire _05604_ ;
wire _05605_ ;
wire _05606_ ;
wire _05607_ ;
wire _05608_ ;
wire _05609_ ;
wire _05610_ ;
wire _05611_ ;
wire _05612_ ;
wire _05613_ ;
wire _05614_ ;
wire _05615_ ;
wire _05616_ ;
wire _05617_ ;
wire _05618_ ;
wire _05619_ ;
wire _05620_ ;
wire _05621_ ;
wire _05622_ ;
wire _05623_ ;
wire _05624_ ;
wire _05625_ ;
wire _05626_ ;
wire _05627_ ;
wire _05628_ ;
wire _05629_ ;
wire _05630_ ;
wire _05631_ ;
wire _05632_ ;
wire _05633_ ;
wire _05634_ ;
wire _05635_ ;
wire _05636_ ;
wire _05637_ ;
wire _05638_ ;
wire _05639_ ;
wire _05640_ ;
wire _05641_ ;
wire _05642_ ;
wire _05643_ ;
wire _05644_ ;
wire _05645_ ;
wire _05646_ ;
wire _05647_ ;
wire _05648_ ;
wire _05649_ ;
wire _05650_ ;
wire _05651_ ;
wire _05652_ ;
wire _05653_ ;
wire _05654_ ;
wire _05655_ ;
wire _05656_ ;
wire _05657_ ;
wire _05658_ ;
wire _05659_ ;
wire _05660_ ;
wire _05661_ ;
wire _05662_ ;
wire _05663_ ;
wire _05664_ ;
wire _05665_ ;
wire _05666_ ;
wire _05667_ ;
wire _05668_ ;
wire _05669_ ;
wire _05670_ ;
wire _05671_ ;
wire _05672_ ;
wire _05673_ ;
wire _05674_ ;
wire _05675_ ;
wire _05676_ ;
wire _05677_ ;
wire _05678_ ;
wire _05679_ ;
wire _05680_ ;
wire _05681_ ;
wire _05682_ ;
wire _05683_ ;
wire _05684_ ;
wire _05685_ ;
wire _05686_ ;
wire _05687_ ;
wire _05688_ ;
wire _05689_ ;
wire _05690_ ;
wire _05691_ ;
wire _05692_ ;
wire _05693_ ;
wire _05694_ ;
wire _05695_ ;
wire _05696_ ;
wire _05697_ ;
wire _05698_ ;
wire _05699_ ;
wire _05700_ ;
wire _05701_ ;
wire _05702_ ;
wire _05703_ ;
wire _05704_ ;
wire _05705_ ;
wire _05706_ ;
wire _05707_ ;
wire _05708_ ;
wire _05709_ ;
wire _05710_ ;
wire _05711_ ;
wire _05712_ ;
wire _05713_ ;
wire _05714_ ;
wire _05715_ ;
wire _05716_ ;
wire _05717_ ;
wire _05718_ ;
wire _05719_ ;
wire _05720_ ;
wire _05721_ ;
wire _05722_ ;
wire _05723_ ;
wire _05724_ ;
wire _05725_ ;
wire _05726_ ;
wire _05727_ ;
wire _05728_ ;
wire _05729_ ;
wire _05730_ ;
wire _05731_ ;
wire _05732_ ;
wire _05733_ ;
wire _05734_ ;
wire _05735_ ;
wire _05736_ ;
wire _05737_ ;
wire _05738_ ;
wire _05739_ ;
wire _05740_ ;
wire _05741_ ;
wire _05742_ ;
wire _05743_ ;
wire _05744_ ;
wire _05745_ ;
wire _05746_ ;
wire _05747_ ;
wire _05748_ ;
wire _05749_ ;
wire _05750_ ;
wire _05751_ ;
wire _05752_ ;
wire _05753_ ;
wire _05754_ ;
wire _05755_ ;
wire _05756_ ;
wire _05757_ ;
wire _05758_ ;
wire _05759_ ;
wire _05760_ ;
wire _05761_ ;
wire _05762_ ;
wire _05763_ ;
wire _05764_ ;
wire _05765_ ;
wire _05766_ ;
wire _05767_ ;
wire _05768_ ;
wire _05769_ ;
wire _05770_ ;
wire _05771_ ;
wire _05772_ ;
wire _05773_ ;
wire _05774_ ;
wire _05775_ ;
wire _05776_ ;
wire _05777_ ;
wire _05778_ ;
wire _05779_ ;
wire _05780_ ;
wire _05781_ ;
wire _05782_ ;
wire _05783_ ;
wire _05784_ ;
wire _05785_ ;
wire _05786_ ;
wire _05787_ ;
wire _05788_ ;
wire _05789_ ;
wire _05790_ ;
wire _05791_ ;
wire _05792_ ;
wire _05793_ ;
wire _05794_ ;
wire _05795_ ;
wire _05796_ ;
wire _05797_ ;
wire _05798_ ;
wire _05799_ ;
wire _05800_ ;
wire _05801_ ;
wire _05802_ ;
wire _05803_ ;
wire _05804_ ;
wire _05805_ ;
wire _05806_ ;
wire _05807_ ;
wire _05808_ ;
wire _05809_ ;
wire _05810_ ;
wire _05811_ ;
wire _05812_ ;
wire _05813_ ;
wire _05814_ ;
wire _05815_ ;
wire _05816_ ;
wire _05817_ ;
wire _05818_ ;
wire _05819_ ;
wire _05820_ ;
wire _05821_ ;
wire _05822_ ;
wire _05823_ ;
wire _05824_ ;
wire _05825_ ;
wire _05826_ ;
wire _05827_ ;
wire _05828_ ;
wire _05829_ ;
wire _05830_ ;
wire _05831_ ;
wire _05832_ ;
wire _05833_ ;
wire _05834_ ;
wire _05835_ ;
wire _05836_ ;
wire _05837_ ;
wire _05838_ ;
wire _05839_ ;
wire _05840_ ;
wire _05841_ ;
wire _05842_ ;
wire _05843_ ;
wire _05844_ ;
wire _05845_ ;
wire _05846_ ;
wire _05847_ ;
wire _05848_ ;
wire _05849_ ;
wire _05850_ ;
wire _05851_ ;
wire _05852_ ;
wire _05853_ ;
wire _05854_ ;
wire _05855_ ;
wire _05856_ ;
wire _05857_ ;
wire _05858_ ;
wire _05859_ ;
wire _05860_ ;
wire _05861_ ;
wire _05862_ ;
wire _05863_ ;
wire _05864_ ;
wire _05865_ ;
wire _05866_ ;
wire _05867_ ;
wire _05868_ ;
wire _05869_ ;
wire _05870_ ;
wire _05871_ ;
wire _05872_ ;
wire _05873_ ;
wire _05874_ ;
wire _05875_ ;
wire _05876_ ;
wire _05877_ ;
wire _05878_ ;
wire _05879_ ;
wire _05880_ ;
wire _05881_ ;
wire _05882_ ;
wire _05883_ ;
wire _05884_ ;
wire _05885_ ;
wire _05886_ ;
wire _05887_ ;
wire _05888_ ;
wire _05889_ ;
wire _05890_ ;
wire _05891_ ;
wire _05892_ ;
wire _05893_ ;
wire _05894_ ;
wire _05895_ ;
wire _05896_ ;
wire _05897_ ;
wire _05898_ ;
wire _05899_ ;
wire _05900_ ;
wire _05901_ ;
wire _05902_ ;
wire _05903_ ;
wire _05904_ ;
wire _05905_ ;
wire _05906_ ;
wire _05907_ ;
wire _05908_ ;
wire _05909_ ;
wire _05910_ ;
wire _05911_ ;
wire _05912_ ;
wire _05913_ ;
wire _05914_ ;
wire _05915_ ;
wire _05916_ ;
wire _05917_ ;
wire _05918_ ;
wire _05919_ ;
wire _05920_ ;
wire _05921_ ;
wire _05922_ ;
wire _05923_ ;
wire _05924_ ;
wire _05925_ ;
wire _05926_ ;
wire _05927_ ;
wire _05928_ ;
wire _05929_ ;
wire _05930_ ;
wire _05931_ ;
wire _05932_ ;
wire _05933_ ;
wire _05934_ ;
wire _05935_ ;
wire _05936_ ;
wire _05937_ ;
wire _05938_ ;
wire _05939_ ;
wire _05940_ ;
wire _05941_ ;
wire _05942_ ;
wire _05943_ ;
wire _05944_ ;
wire _05945_ ;
wire _05946_ ;
wire _05947_ ;
wire _05948_ ;
wire _05949_ ;
wire _05950_ ;
wire _05951_ ;
wire _05952_ ;
wire _05953_ ;
wire _05954_ ;
wire _05955_ ;
wire _05956_ ;
wire _05957_ ;
wire _05958_ ;
wire _05959_ ;
wire _05960_ ;
wire _05961_ ;
wire _05962_ ;
wire _05963_ ;
wire _05964_ ;
wire _05965_ ;
wire _05966_ ;
wire _05967_ ;
wire _05968_ ;
wire _05969_ ;
wire _05970_ ;
wire _05971_ ;
wire _05972_ ;
wire _05973_ ;
wire _05974_ ;
wire _05975_ ;
wire _05976_ ;
wire _05977_ ;
wire _05978_ ;
wire _05979_ ;
wire _05980_ ;
wire _05981_ ;
wire _05982_ ;
wire _05983_ ;
wire _05984_ ;
wire _05985_ ;
wire _05986_ ;
wire _05987_ ;
wire _05988_ ;
wire _05989_ ;
wire _05990_ ;
wire _05991_ ;
wire _05992_ ;
wire _05993_ ;
wire _05994_ ;
wire _05995_ ;
wire _05996_ ;
wire _05997_ ;
wire _05998_ ;
wire _05999_ ;
wire _06000_ ;
wire _06001_ ;
wire _06002_ ;
wire _06003_ ;
wire _06004_ ;
wire _06005_ ;
wire _06006_ ;
wire _06007_ ;
wire _06008_ ;
wire _06009_ ;
wire _06010_ ;
wire _06011_ ;
wire _06012_ ;
wire _06013_ ;
wire _06014_ ;
wire _06015_ ;
wire _06016_ ;
wire _06017_ ;
wire _06018_ ;
wire _06019_ ;
wire _06020_ ;
wire _06021_ ;
wire _06022_ ;
wire _06023_ ;
wire _06024_ ;
wire _06025_ ;
wire _06026_ ;
wire _06027_ ;
wire _06028_ ;
wire _06029_ ;
wire _06030_ ;
wire _06031_ ;
wire _06032_ ;
wire _06033_ ;
wire _06034_ ;
wire _06035_ ;
wire _06036_ ;
wire _06037_ ;
wire _06038_ ;
wire _06039_ ;
wire _06040_ ;
wire _06041_ ;
wire _06042_ ;
wire _06043_ ;
wire _06044_ ;
wire _06045_ ;
wire _06046_ ;
wire _06047_ ;
wire _06048_ ;
wire _06049_ ;
wire _06050_ ;
wire _06051_ ;
wire _06052_ ;
wire _06053_ ;
wire _06054_ ;
wire _06055_ ;
wire _06056_ ;
wire _06057_ ;
wire _06058_ ;
wire _06059_ ;
wire _06060_ ;
wire _06061_ ;
wire _06062_ ;
wire _06063_ ;
wire _06064_ ;
wire _06065_ ;
wire _06066_ ;
wire _06067_ ;
wire _06068_ ;
wire _06069_ ;
wire _06070_ ;
wire _06071_ ;
wire _06072_ ;
wire _06073_ ;
wire _06074_ ;
wire _06075_ ;
wire _06076_ ;
wire _06077_ ;
wire _06078_ ;
wire _06079_ ;
wire _06080_ ;
wire _06081_ ;
wire _06082_ ;
wire _06083_ ;
wire _06084_ ;
wire _06085_ ;
wire _06086_ ;
wire _06087_ ;
wire _06088_ ;
wire _06089_ ;
wire _06090_ ;
wire _06091_ ;
wire _06092_ ;
wire _06093_ ;
wire _06094_ ;
wire _06095_ ;
wire _06096_ ;
wire _06097_ ;
wire _06098_ ;
wire _06099_ ;
wire _06100_ ;
wire _06101_ ;
wire _06102_ ;
wire _06103_ ;
wire _06104_ ;
wire _06105_ ;
wire _06106_ ;
wire _06107_ ;
wire _06108_ ;
wire _06109_ ;
wire _06110_ ;
wire _06111_ ;
wire _06112_ ;
wire _06113_ ;
wire _06114_ ;
wire _06115_ ;
wire _06116_ ;
wire _06117_ ;
wire _06118_ ;
wire _06119_ ;
wire _06120_ ;
wire _06121_ ;
wire _06122_ ;
wire _06123_ ;
wire _06124_ ;
wire _06125_ ;
wire _06126_ ;
wire _06127_ ;
wire _06128_ ;
wire _06129_ ;
wire _06130_ ;
wire _06131_ ;
wire _06132_ ;
wire _06133_ ;
wire _06134_ ;
wire _06135_ ;
wire _06136_ ;
wire _06137_ ;
wire _06138_ ;
wire _06139_ ;
wire _06140_ ;
wire _06141_ ;
wire _06142_ ;
wire _06143_ ;
wire _06144_ ;
wire _06145_ ;
wire _06146_ ;
wire _06147_ ;
wire _06148_ ;
wire _06149_ ;
wire _06150_ ;
wire _06151_ ;
wire _06152_ ;
wire _06153_ ;
wire _06154_ ;
wire _06155_ ;
wire _06156_ ;
wire _06157_ ;
wire _06158_ ;
wire _06159_ ;
wire _06160_ ;
wire _06161_ ;
wire _06162_ ;
wire _06163_ ;
wire _06164_ ;
wire _06165_ ;
wire _06166_ ;
wire _06167_ ;
wire _06168_ ;
wire _06169_ ;
wire _06170_ ;
wire _06171_ ;
wire _06172_ ;
wire _06173_ ;
wire _06174_ ;
wire _06175_ ;
wire _06176_ ;
wire _06177_ ;
wire _06178_ ;
wire _06179_ ;
wire _06180_ ;
wire _06181_ ;
wire _06182_ ;
wire _06183_ ;
wire _06184_ ;
wire _06185_ ;
wire _06186_ ;
wire _06187_ ;
wire _06188_ ;
wire _06189_ ;
wire _06190_ ;
wire _06191_ ;
wire _06192_ ;
wire _06193_ ;
wire _06194_ ;
wire _06195_ ;
wire _06196_ ;
wire _06197_ ;
wire _06198_ ;
wire _06199_ ;
wire _06200_ ;
wire _06201_ ;
wire _06202_ ;
wire _06203_ ;
wire _06204_ ;
wire _06205_ ;
wire _06206_ ;
wire _06207_ ;
wire _06208_ ;
wire _06209_ ;
wire _06210_ ;
wire _06211_ ;
wire _06212_ ;
wire _06213_ ;
wire _06214_ ;
wire _06215_ ;
wire _06216_ ;
wire _06217_ ;
wire _06218_ ;
wire _06219_ ;
wire _06220_ ;
wire _06221_ ;
wire _06222_ ;
wire _06223_ ;
wire _06224_ ;
wire _06225_ ;
wire _06226_ ;
wire _06227_ ;
wire _06228_ ;
wire _06229_ ;
wire _06230_ ;
wire _06231_ ;
wire _06232_ ;
wire _06233_ ;
wire _06234_ ;
wire _06235_ ;
wire _06236_ ;
wire _06237_ ;
wire _06238_ ;
wire _06239_ ;
wire _06240_ ;
wire _06241_ ;
wire _06242_ ;
wire _06243_ ;
wire _06244_ ;
wire _06245_ ;
wire _06246_ ;
wire _06247_ ;
wire _06248_ ;
wire _06249_ ;
wire _06250_ ;
wire _06251_ ;
wire _06252_ ;
wire _06253_ ;
wire _06254_ ;
wire _06255_ ;
wire _06256_ ;
wire _06257_ ;
wire _06258_ ;
wire _06259_ ;
wire _06260_ ;
wire _06261_ ;
wire _06262_ ;
wire _06263_ ;
wire _06264_ ;
wire _06265_ ;
wire _06266_ ;
wire _06267_ ;
wire _06268_ ;
wire _06269_ ;
wire _06270_ ;
wire _06271_ ;
wire _06272_ ;
wire _06273_ ;
wire _06274_ ;
wire _06275_ ;
wire _06276_ ;
wire _06277_ ;
wire _06278_ ;
wire _06279_ ;
wire _06280_ ;
wire _06281_ ;
wire _06282_ ;
wire _06283_ ;
wire _06284_ ;
wire _06285_ ;
wire _06286_ ;
wire _06287_ ;
wire _06288_ ;
wire _06289_ ;
wire _06290_ ;
wire _06291_ ;
wire _06292_ ;
wire _06293_ ;
wire _06294_ ;
wire _06295_ ;
wire _06296_ ;
wire _06297_ ;
wire _06298_ ;
wire _06299_ ;
wire _06300_ ;
wire _06301_ ;
wire _06302_ ;
wire _06303_ ;
wire _06304_ ;
wire _06305_ ;
wire _06306_ ;
wire _06307_ ;
wire _06308_ ;
wire _06309_ ;
wire _06310_ ;
wire _06311_ ;
wire _06312_ ;
wire _06313_ ;
wire _06314_ ;
wire _06315_ ;
wire _06316_ ;
wire _06317_ ;
wire _06318_ ;
wire _06319_ ;
wire _06320_ ;
wire _06321_ ;
wire _06322_ ;
wire _06323_ ;
wire _06324_ ;
wire _06325_ ;
wire _06326_ ;
wire _06327_ ;
wire _06328_ ;
wire _06329_ ;
wire _06330_ ;
wire _06331_ ;
wire _06332_ ;
wire _06333_ ;
wire _06334_ ;
wire _06335_ ;
wire _06336_ ;
wire _06337_ ;
wire _06338_ ;
wire _06339_ ;
wire _06340_ ;
wire _06341_ ;
wire _06342_ ;
wire _06343_ ;
wire _06344_ ;
wire _06345_ ;
wire _06346_ ;
wire _06347_ ;
wire _06348_ ;
wire _06349_ ;
wire _06350_ ;
wire _06351_ ;
wire _06352_ ;
wire _06353_ ;
wire _06354_ ;
wire _06355_ ;
wire _06356_ ;
wire _06357_ ;
wire _06358_ ;
wire _06359_ ;
wire _06360_ ;
wire _06361_ ;
wire _06362_ ;
wire _06363_ ;
wire _06364_ ;
wire _06365_ ;
wire _06366_ ;
wire _06367_ ;
wire _06368_ ;
wire _06369_ ;
wire _06370_ ;
wire _06371_ ;
wire _06372_ ;
wire _06373_ ;
wire _06374_ ;
wire _06375_ ;
wire _06376_ ;
wire _06377_ ;
wire _06378_ ;
wire _06379_ ;
wire _06380_ ;
wire _06381_ ;
wire _06382_ ;
wire _06383_ ;
wire _06384_ ;
wire _06385_ ;
wire _06386_ ;
wire _06387_ ;
wire _06388_ ;
wire _06389_ ;
wire _06390_ ;
wire _06391_ ;
wire _06392_ ;
wire _06393_ ;
wire _06394_ ;
wire _06395_ ;
wire _06396_ ;
wire _06397_ ;
wire _06398_ ;
wire _06399_ ;
wire _06400_ ;
wire _06401_ ;
wire _06402_ ;
wire _06403_ ;
wire _06404_ ;
wire _06405_ ;
wire _06406_ ;
wire _06407_ ;
wire _06408_ ;
wire _06409_ ;
wire _06410_ ;
wire _06411_ ;
wire _06412_ ;
wire _06413_ ;
wire _06414_ ;
wire _06415_ ;
wire _06416_ ;
wire _06417_ ;
wire _06418_ ;
wire _06419_ ;
wire _06420_ ;
wire _06421_ ;
wire _06422_ ;
wire _06423_ ;
wire _06424_ ;
wire _06425_ ;
wire _06426_ ;
wire _06427_ ;
wire _06428_ ;
wire _06429_ ;
wire _06430_ ;
wire _06431_ ;
wire _06432_ ;
wire _06433_ ;
wire _06434_ ;
wire _06435_ ;
wire _06436_ ;
wire _06437_ ;
wire _06438_ ;
wire _06439_ ;
wire _06440_ ;
wire _06441_ ;
wire _06442_ ;
wire _06443_ ;
wire _06444_ ;
wire _06445_ ;
wire _06446_ ;
wire _06447_ ;
wire _06448_ ;
wire _06449_ ;
wire _06450_ ;
wire _06451_ ;
wire _06452_ ;
wire _06453_ ;
wire _06454_ ;
wire _06455_ ;
wire _06456_ ;
wire _06457_ ;
wire _06458_ ;
wire _06459_ ;
wire _06460_ ;
wire _06461_ ;
wire _06462_ ;
wire _06463_ ;
wire _06464_ ;
wire _06465_ ;
wire _06466_ ;
wire _06467_ ;
wire _06468_ ;
wire _06469_ ;
wire _06470_ ;
wire _06471_ ;
wire _06472_ ;
wire _06473_ ;
wire _06474_ ;
wire _06475_ ;
wire _06476_ ;
wire _06477_ ;
wire _06478_ ;
wire _06479_ ;
wire _06480_ ;
wire _06481_ ;
wire _06482_ ;
wire _06483_ ;
wire _06484_ ;
wire _06485_ ;
wire _06486_ ;
wire _06487_ ;
wire _06488_ ;
wire _06489_ ;
wire _06490_ ;
wire _06491_ ;
wire _06492_ ;
wire _06493_ ;
wire _06494_ ;
wire _06495_ ;
wire _06496_ ;
wire _06497_ ;
wire _06498_ ;
wire _06499_ ;
wire _06500_ ;
wire _06501_ ;
wire _06502_ ;
wire _06503_ ;
wire _06504_ ;
wire _06505_ ;
wire _06506_ ;
wire _06507_ ;
wire _06508_ ;
wire _06509_ ;
wire _06510_ ;
wire _06511_ ;
wire _06512_ ;
wire _06513_ ;
wire _06514_ ;
wire _06515_ ;
wire _06516_ ;
wire _06517_ ;
wire _06518_ ;
wire _06519_ ;
wire _06520_ ;
wire _06521_ ;
wire _06522_ ;
wire _06523_ ;
wire _06524_ ;
wire _06525_ ;
wire _06526_ ;
wire _06527_ ;
wire _06528_ ;
wire _06529_ ;
wire _06530_ ;
wire _06531_ ;
wire _06532_ ;
wire _06533_ ;
wire _06534_ ;
wire _06535_ ;
wire _06536_ ;
wire _06537_ ;
wire _06538_ ;
wire _06539_ ;
wire _06540_ ;
wire _06541_ ;
wire _06542_ ;
wire _06543_ ;
wire _06544_ ;
wire _06545_ ;
wire _06546_ ;
wire _06547_ ;
wire _06548_ ;
wire _06549_ ;
wire _06550_ ;
wire _06551_ ;
wire _06552_ ;
wire _06553_ ;
wire _06554_ ;
wire _06555_ ;
wire _06556_ ;
wire _06557_ ;
wire _06558_ ;
wire _06559_ ;
wire _06560_ ;
wire _06561_ ;
wire _06562_ ;
wire _06563_ ;
wire _06564_ ;
wire _06565_ ;
wire _06566_ ;
wire _06567_ ;
wire _06568_ ;
wire _06569_ ;
wire _06570_ ;
wire _06571_ ;
wire _06572_ ;
wire _06573_ ;
wire _06574_ ;
wire _06575_ ;
wire _06576_ ;
wire _06577_ ;
wire _06578_ ;
wire _06579_ ;
wire _06580_ ;
wire _06581_ ;
wire _06582_ ;
wire _06583_ ;
wire _06584_ ;
wire _06585_ ;
wire _06586_ ;
wire _06587_ ;
wire _06588_ ;
wire _06589_ ;
wire _06590_ ;
wire _06591_ ;
wire _06592_ ;
wire _06593_ ;
wire _06594_ ;
wire _06595_ ;
wire _06596_ ;
wire _06597_ ;
wire _06598_ ;
wire _06599_ ;
wire _06600_ ;
wire _06601_ ;
wire _06602_ ;
wire _06603_ ;
wire _06604_ ;
wire _06605_ ;
wire _06606_ ;
wire _06607_ ;
wire _06608_ ;
wire _06609_ ;
wire _06610_ ;
wire _06611_ ;
wire _06612_ ;
wire _06613_ ;
wire _06614_ ;
wire _06615_ ;
wire _06616_ ;
wire _06617_ ;
wire _06618_ ;
wire _06619_ ;
wire _06620_ ;
wire _06621_ ;
wire _06622_ ;
wire _06623_ ;
wire _06624_ ;
wire _06625_ ;
wire _06626_ ;
wire _06627_ ;
wire _06628_ ;
wire _06629_ ;
wire _06630_ ;
wire _06631_ ;
wire _06632_ ;
wire _06633_ ;
wire _06634_ ;
wire _06635_ ;
wire _06636_ ;
wire _06637_ ;
wire _06638_ ;
wire _06639_ ;
wire _06640_ ;
wire _06641_ ;
wire _06642_ ;
wire _06643_ ;
wire _06644_ ;
wire _06645_ ;
wire _06646_ ;
wire _06647_ ;
wire _06648_ ;
wire _06649_ ;
wire _06650_ ;
wire _06651_ ;
wire _06652_ ;
wire _06653_ ;
wire _06654_ ;
wire _06655_ ;
wire _06656_ ;
wire _06657_ ;
wire _06658_ ;
wire _06659_ ;
wire _06660_ ;
wire _06661_ ;
wire _06662_ ;
wire _06663_ ;
wire _06664_ ;
wire _06665_ ;
wire _06666_ ;
wire _06667_ ;
wire _06668_ ;
wire _06669_ ;
wire _06670_ ;
wire _06671_ ;
wire _06672_ ;
wire _06673_ ;
wire _06674_ ;
wire _06675_ ;
wire _06676_ ;
wire _06677_ ;
wire _06678_ ;
wire _06679_ ;
wire _06680_ ;
wire _06681_ ;
wire _06682_ ;
wire _06683_ ;
wire _06684_ ;
wire _06685_ ;
wire _06686_ ;
wire _06687_ ;
wire _06688_ ;
wire _06689_ ;
wire _06690_ ;
wire _06691_ ;
wire _06692_ ;
wire _06693_ ;
wire _06694_ ;
wire _06695_ ;
wire _06696_ ;
wire _06697_ ;
wire _06698_ ;
wire _06699_ ;
wire _06700_ ;
wire _06701_ ;
wire _06702_ ;
wire _06703_ ;
wire _06704_ ;
wire _06705_ ;
wire _06706_ ;
wire _06707_ ;
wire _06708_ ;
wire _06709_ ;
wire _06710_ ;
wire _06711_ ;
wire _06712_ ;
wire _06713_ ;
wire _06714_ ;
wire _06715_ ;
wire _06716_ ;
wire _06717_ ;
wire _06718_ ;
wire _06719_ ;
wire _06720_ ;
wire _06721_ ;
wire _06722_ ;
wire _06723_ ;
wire _06724_ ;
wire _06725_ ;
wire _06726_ ;
wire _06727_ ;
wire _06728_ ;
wire _06729_ ;
wire _06730_ ;
wire _06731_ ;
wire _06732_ ;
wire _06733_ ;
wire _06734_ ;
wire _06735_ ;
wire _06736_ ;
wire _06737_ ;
wire _06738_ ;
wire _06739_ ;
wire _06740_ ;
wire _06741_ ;
wire _06742_ ;
wire _06743_ ;
wire _06744_ ;
wire _06745_ ;
wire _06746_ ;
wire _06747_ ;
wire _06748_ ;
wire _06749_ ;
wire _06750_ ;
wire _06751_ ;
wire _06752_ ;
wire _06753_ ;
wire _06754_ ;
wire _06755_ ;
wire _06756_ ;
wire _06757_ ;
wire _06758_ ;
wire _06759_ ;
wire _06760_ ;
wire _06761_ ;
wire _06762_ ;
wire _06763_ ;
wire _06764_ ;
wire _06765_ ;
wire _06766_ ;
wire _06767_ ;
wire _06768_ ;
wire _06769_ ;
wire _06770_ ;
wire _06771_ ;
wire _06772_ ;
wire _06773_ ;
wire _06774_ ;
wire _06775_ ;
wire _06776_ ;
wire _06777_ ;
wire _06778_ ;
wire _06779_ ;
wire _06780_ ;
wire _06781_ ;
wire _06782_ ;
wire _06783_ ;
wire _06784_ ;
wire _06785_ ;
wire _06786_ ;
wire _06787_ ;
wire _06788_ ;
wire _06789_ ;
wire _06790_ ;
wire _06791_ ;
wire _06792_ ;
wire _06793_ ;
wire _06794_ ;
wire _06795_ ;
wire _06796_ ;
wire _06797_ ;
wire _06798_ ;
wire _06799_ ;
wire _06800_ ;
wire _06801_ ;
wire _06802_ ;
wire _06803_ ;
wire _06804_ ;
wire _06805_ ;
wire _06806_ ;
wire _06807_ ;
wire _06808_ ;
wire _06809_ ;
wire _06810_ ;
wire _06811_ ;
wire _06812_ ;
wire _06813_ ;
wire _06814_ ;
wire _06815_ ;
wire _06816_ ;
wire _06817_ ;
wire _06818_ ;
wire _06819_ ;
wire _06820_ ;
wire _06821_ ;
wire _06822_ ;
wire _06823_ ;
wire _06824_ ;
wire _06825_ ;
wire _06826_ ;
wire _06827_ ;
wire _06828_ ;
wire _06829_ ;
wire _06830_ ;
wire _06831_ ;
wire _06832_ ;
wire _06833_ ;
wire _06834_ ;
wire _06835_ ;
wire _06836_ ;
wire _06837_ ;
wire _06838_ ;
wire _06839_ ;
wire _06840_ ;
wire _06841_ ;
wire _06842_ ;
wire _06843_ ;
wire _06844_ ;
wire _06845_ ;
wire _06846_ ;
wire _06847_ ;
wire _06848_ ;
wire _06849_ ;
wire _06850_ ;
wire _06851_ ;
wire _06852_ ;
wire _06853_ ;
wire _06854_ ;
wire _06855_ ;
wire _06856_ ;
wire _06857_ ;
wire _06858_ ;
wire _06859_ ;
wire _06860_ ;
wire _06861_ ;
wire _06862_ ;
wire _06863_ ;
wire _06864_ ;
wire _06865_ ;
wire _06866_ ;
wire _06867_ ;
wire _06868_ ;
wire _06869_ ;
wire _06870_ ;
wire _06871_ ;
wire _06872_ ;
wire _06873_ ;
wire _06874_ ;
wire _06875_ ;
wire _06876_ ;
wire _06877_ ;
wire _06878_ ;
wire _06879_ ;
wire _06880_ ;
wire _06881_ ;
wire _06882_ ;
wire _06883_ ;
wire _06884_ ;
wire _06885_ ;
wire _06886_ ;
wire _06887_ ;
wire _06888_ ;
wire _06889_ ;
wire _06890_ ;
wire _06891_ ;
wire _06892_ ;
wire _06893_ ;
wire _06894_ ;
wire _06895_ ;
wire _06896_ ;
wire _06897_ ;
wire _06898_ ;
wire _06899_ ;
wire _06900_ ;
wire _06901_ ;
wire _06902_ ;
wire _06903_ ;
wire _06904_ ;
wire _06905_ ;
wire _06906_ ;
wire _06907_ ;
wire _06908_ ;
wire _06909_ ;
wire _06910_ ;
wire _06911_ ;
wire _06912_ ;
wire _06913_ ;
wire _06914_ ;
wire _06915_ ;
wire _06916_ ;
wire _06917_ ;
wire _06918_ ;
wire _06919_ ;
wire _06920_ ;
wire _06921_ ;
wire _06922_ ;
wire _06923_ ;
wire _06924_ ;
wire _06925_ ;
wire _06926_ ;
wire _06927_ ;
wire _06928_ ;
wire _06929_ ;
wire _06930_ ;
wire _06931_ ;
wire _06932_ ;
wire _06933_ ;
wire _06934_ ;
wire _06935_ ;
wire _06936_ ;
wire _06937_ ;
wire _06938_ ;
wire _06939_ ;
wire _06940_ ;
wire _06941_ ;
wire _06942_ ;
wire _06943_ ;
wire _06944_ ;
wire _06945_ ;
wire _06946_ ;
wire _06947_ ;
wire _06948_ ;
wire _06949_ ;
wire _06950_ ;
wire _06951_ ;
wire _06952_ ;
wire _06953_ ;
wire _06954_ ;
wire _06955_ ;
wire _06956_ ;
wire _06957_ ;
wire _06958_ ;
wire _06959_ ;
wire _06960_ ;
wire _06961_ ;
wire _06962_ ;
wire _06963_ ;
wire _06964_ ;
wire _06965_ ;
wire _06966_ ;
wire _06967_ ;
wire _06968_ ;
wire _06969_ ;
wire _06970_ ;
wire _06971_ ;
wire _06972_ ;
wire _06973_ ;
wire _06974_ ;
wire _06975_ ;
wire _06976_ ;
wire _06977_ ;
wire _06978_ ;
wire _06979_ ;
wire _06980_ ;
wire _06981_ ;
wire _06982_ ;
wire _06983_ ;
wire _06984_ ;
wire _06985_ ;
wire _06986_ ;
wire _06987_ ;
wire _06988_ ;
wire _06989_ ;
wire _06990_ ;
wire _06991_ ;
wire _06992_ ;
wire _06993_ ;
wire _06994_ ;
wire _06995_ ;
wire _06996_ ;
wire _06997_ ;
wire _06998_ ;
wire _06999_ ;
wire _07000_ ;
wire _07001_ ;
wire _07002_ ;
wire _07003_ ;
wire _07004_ ;
wire _07005_ ;
wire _07006_ ;
wire _07007_ ;
wire _07008_ ;
wire _07009_ ;
wire _07010_ ;
wire _07011_ ;
wire _07012_ ;
wire _07013_ ;
wire _07014_ ;
wire _07015_ ;
wire _07016_ ;
wire _07017_ ;
wire _07018_ ;
wire _07019_ ;
wire _07020_ ;
wire _07021_ ;
wire _07022_ ;
wire _07023_ ;
wire _07024_ ;
wire _07025_ ;
wire _07026_ ;
wire _07027_ ;
wire _07028_ ;
wire _07029_ ;
wire _07030_ ;
wire _07031_ ;
wire _07032_ ;
wire _07033_ ;
wire _07034_ ;
wire _07035_ ;
wire _07036_ ;
wire _07037_ ;
wire _07038_ ;
wire _07039_ ;
wire _07040_ ;
wire _07041_ ;
wire _07042_ ;
wire _07043_ ;
wire _07044_ ;
wire _07045_ ;
wire _07046_ ;
wire _07047_ ;
wire _07048_ ;
wire _07049_ ;
wire _07050_ ;
wire _07051_ ;
wire _07052_ ;
wire _07053_ ;
wire _07054_ ;
wire _07055_ ;
wire _07056_ ;
wire _07057_ ;
wire _07058_ ;
wire _07059_ ;
wire _07060_ ;
wire _07061_ ;
wire _07062_ ;
wire _07063_ ;
wire _07064_ ;
wire _07065_ ;
wire _07066_ ;
wire _07067_ ;
wire _07068_ ;
wire _07069_ ;
wire _07070_ ;
wire _07071_ ;
wire _07072_ ;
wire _07073_ ;
wire _07074_ ;
wire _07075_ ;
wire _07076_ ;
wire _07077_ ;
wire _07078_ ;
wire _07079_ ;
wire _07080_ ;
wire _07081_ ;
wire _07082_ ;
wire _07083_ ;
wire _07084_ ;
wire _07085_ ;
wire _07086_ ;
wire _07087_ ;
wire _07088_ ;
wire _07089_ ;
wire _07090_ ;
wire _07091_ ;
wire _07092_ ;
wire _07093_ ;
wire _07094_ ;
wire _07095_ ;
wire _07096_ ;
wire _07097_ ;
wire _07098_ ;
wire _07099_ ;
wire _07100_ ;
wire _07101_ ;
wire _07102_ ;
wire _07103_ ;
wire _07104_ ;
wire _07105_ ;
wire _07106_ ;
wire _07107_ ;
wire _07108_ ;
wire _07109_ ;
wire _07110_ ;
wire _07111_ ;
wire _07112_ ;
wire _07113_ ;
wire _07114_ ;
wire _07115_ ;
wire _07116_ ;
wire _07117_ ;
wire _07118_ ;
wire _07119_ ;
wire _07120_ ;
wire _07121_ ;
wire _07122_ ;
wire _07123_ ;
wire _07124_ ;
wire _07125_ ;
wire _07126_ ;
wire _07127_ ;
wire _07128_ ;
wire _07129_ ;
wire _07130_ ;
wire _07131_ ;
wire _07132_ ;
wire _07133_ ;
wire _07134_ ;
wire _07135_ ;
wire _07136_ ;
wire _07137_ ;
wire _07138_ ;
wire _07139_ ;
wire _07140_ ;
wire _07141_ ;
wire _07142_ ;
wire _07143_ ;
wire _07144_ ;
wire _07145_ ;
wire _07146_ ;
wire _07147_ ;
wire _07148_ ;
wire _07149_ ;
wire _07150_ ;
wire _07151_ ;
wire _07152_ ;
wire _07153_ ;
wire _07154_ ;
wire _07155_ ;
wire _07156_ ;
wire _07157_ ;
wire _07158_ ;
wire _07159_ ;
wire _07160_ ;
wire _07161_ ;
wire _07162_ ;
wire _07163_ ;
wire _07164_ ;
wire _07165_ ;
wire _07166_ ;
wire _07167_ ;
wire _07168_ ;
wire _07169_ ;
wire _07170_ ;
wire _07171_ ;
wire _07172_ ;
wire _07173_ ;
wire _07174_ ;
wire _07175_ ;
wire _07176_ ;
wire _07177_ ;
wire _07178_ ;
wire _07179_ ;
wire _07180_ ;
wire _07181_ ;
wire _07182_ ;
wire _07183_ ;
wire _07184_ ;
wire _07185_ ;
wire _07186_ ;
wire _07187_ ;
wire _07188_ ;
wire _07189_ ;
wire _07190_ ;
wire _07191_ ;
wire _07192_ ;
wire _07193_ ;
wire _07194_ ;
wire _07195_ ;
wire _07196_ ;
wire _07197_ ;
wire _07198_ ;
wire _07199_ ;
wire _07200_ ;
wire _07201_ ;
wire _07202_ ;
wire _07203_ ;
wire _07204_ ;
wire _07205_ ;
wire _07206_ ;
wire _07207_ ;
wire _07208_ ;
wire _07209_ ;
wire _07210_ ;
wire _07211_ ;
wire _07212_ ;
wire _07213_ ;
wire _07214_ ;
wire _07215_ ;
wire _07216_ ;
wire _07217_ ;
wire _07218_ ;
wire _07219_ ;
wire _07220_ ;
wire _07221_ ;
wire _07222_ ;
wire _07223_ ;
wire _07224_ ;
wire _07225_ ;
wire _07226_ ;
wire _07227_ ;
wire _07228_ ;
wire _07229_ ;
wire _07230_ ;
wire _07231_ ;
wire _07232_ ;
wire _07233_ ;
wire _07234_ ;
wire _07235_ ;
wire _07236_ ;
wire _07237_ ;
wire _07238_ ;
wire _07239_ ;
wire _07240_ ;
wire _07241_ ;
wire _07242_ ;
wire _07243_ ;
wire _07244_ ;
wire _07245_ ;
wire _07246_ ;
wire _07247_ ;
wire _07248_ ;
wire _07249_ ;
wire _07250_ ;
wire _07251_ ;
wire _07252_ ;
wire _07253_ ;
wire _07254_ ;
wire _07255_ ;
wire _07256_ ;
wire _07257_ ;
wire _07258_ ;
wire _07259_ ;
wire _07260_ ;
wire _07261_ ;
wire _07262_ ;
wire _07263_ ;
wire _07264_ ;
wire _07265_ ;
wire _07266_ ;
wire _07267_ ;
wire _07268_ ;
wire _07269_ ;
wire _07270_ ;
wire _07271_ ;
wire _07272_ ;
wire _07273_ ;
wire _07274_ ;
wire _07275_ ;
wire _07276_ ;
wire _07277_ ;
wire _07278_ ;
wire _07279_ ;
wire _07280_ ;
wire _07281_ ;
wire _07282_ ;
wire _07283_ ;
wire _07284_ ;
wire _07285_ ;
wire _07286_ ;
wire _07287_ ;
wire _07288_ ;
wire _07289_ ;
wire _07290_ ;
wire _07291_ ;
wire _07292_ ;
wire _07293_ ;
wire _07294_ ;
wire _07295_ ;
wire _07296_ ;
wire _07297_ ;
wire _07298_ ;
wire _07299_ ;
wire _07300_ ;
wire _07301_ ;
wire _07302_ ;
wire _07303_ ;
wire _07304_ ;
wire _07305_ ;
wire _07306_ ;
wire _07307_ ;
wire _07308_ ;
wire _07309_ ;
wire _07310_ ;
wire _07311_ ;
wire _07312_ ;
wire _07313_ ;
wire _07314_ ;
wire _07315_ ;
wire _07316_ ;
wire _07317_ ;
wire _07318_ ;
wire _07319_ ;
wire _07320_ ;
wire _07321_ ;
wire _07322_ ;
wire _07323_ ;
wire _07324_ ;
wire _07325_ ;
wire _07326_ ;
wire _07327_ ;
wire _07328_ ;
wire _07329_ ;
wire _07330_ ;
wire _07331_ ;
wire _07332_ ;
wire _07333_ ;
wire _07334_ ;
wire _07335_ ;
wire _07336_ ;
wire _07337_ ;
wire _07338_ ;
wire _07339_ ;
wire _07340_ ;
wire _07341_ ;
wire _07342_ ;
wire _07343_ ;
wire _07344_ ;
wire _07345_ ;
wire _07346_ ;
wire _07347_ ;
wire _07348_ ;
wire _07349_ ;
wire _07350_ ;
wire _07351_ ;
wire _07352_ ;
wire _07353_ ;
wire _07354_ ;
wire _07355_ ;
wire _07356_ ;
wire _07357_ ;
wire _07358_ ;
wire _07359_ ;
wire _07360_ ;
wire _07361_ ;
wire _07362_ ;
wire _07363_ ;
wire _07364_ ;
wire _07365_ ;
wire _07366_ ;
wire _07367_ ;
wire _07368_ ;
wire _07369_ ;
wire _07370_ ;
wire _07371_ ;
wire _07372_ ;
wire _07373_ ;
wire _07374_ ;
wire _07375_ ;
wire _07376_ ;
wire _07377_ ;
wire _07378_ ;
wire _07379_ ;
wire _07380_ ;
wire _07381_ ;
wire _07382_ ;
wire _07383_ ;
wire _07384_ ;
wire _07385_ ;
wire _07386_ ;
wire _07387_ ;
wire _07388_ ;
wire _07389_ ;
wire _07390_ ;
wire _07391_ ;
wire _07392_ ;
wire _07393_ ;
wire _07394_ ;
wire _07395_ ;
wire _07396_ ;
wire _07397_ ;
wire _07398_ ;
wire _07399_ ;
wire _07400_ ;
wire _07401_ ;
wire _07402_ ;
wire _07403_ ;
wire _07404_ ;
wire _07405_ ;
wire _07406_ ;
wire _07407_ ;
wire _07408_ ;
wire _07409_ ;
wire _07410_ ;
wire _07411_ ;
wire _07412_ ;
wire _07413_ ;
wire _07414_ ;
wire _07415_ ;
wire _07416_ ;
wire _07417_ ;
wire _07418_ ;
wire _07419_ ;
wire _07420_ ;
wire _07421_ ;
wire _07422_ ;
wire _07423_ ;
wire _07424_ ;
wire _07425_ ;
wire _07426_ ;
wire _07427_ ;
wire _07428_ ;
wire _07429_ ;
wire _07430_ ;
wire _07431_ ;
wire _07432_ ;
wire _07433_ ;
wire _07434_ ;
wire _07435_ ;
wire _07436_ ;
wire _07437_ ;
wire _07438_ ;
wire _07439_ ;
wire _07440_ ;
wire _07441_ ;
wire _07442_ ;
wire _07443_ ;
wire _07444_ ;
wire _07445_ ;
wire _07446_ ;
wire _07447_ ;
wire _07448_ ;
wire _07449_ ;
wire _07450_ ;
wire _07451_ ;
wire _07452_ ;
wire _07453_ ;
wire _07454_ ;
wire _07455_ ;
wire _07456_ ;
wire _07457_ ;
wire _07458_ ;
wire _07459_ ;
wire _07460_ ;
wire _07461_ ;
wire _07462_ ;
wire _07463_ ;
wire _07464_ ;
wire _07465_ ;
wire _07466_ ;
wire _07467_ ;
wire _07468_ ;
wire _07469_ ;
wire _07470_ ;
wire _07471_ ;
wire _07472_ ;
wire _07473_ ;
wire _07474_ ;
wire _07475_ ;
wire _07476_ ;
wire _07477_ ;
wire _07478_ ;
wire _07479_ ;
wire _07480_ ;
wire _07481_ ;
wire _07482_ ;
wire _07483_ ;
wire _07484_ ;
wire _07485_ ;
wire _07486_ ;
wire _07487_ ;
wire _07488_ ;
wire _07489_ ;
wire _07490_ ;
wire _07491_ ;
wire _07492_ ;
wire _07493_ ;
wire _07494_ ;
wire _07495_ ;
wire _07496_ ;
wire _07497_ ;
wire _07498_ ;
wire _07499_ ;
wire _07500_ ;
wire _07501_ ;
wire _07502_ ;
wire _07503_ ;
wire _07504_ ;
wire _07505_ ;
wire _07506_ ;
wire _07507_ ;
wire _07508_ ;
wire _07509_ ;
wire _07510_ ;
wire _07511_ ;
wire _07512_ ;
wire _07513_ ;
wire _07514_ ;
wire _07515_ ;
wire _07516_ ;
wire _07517_ ;
wire _07518_ ;
wire _07519_ ;
wire _07520_ ;
wire _07521_ ;
wire _07522_ ;
wire _07523_ ;
wire _07524_ ;
wire _07525_ ;
wire _07526_ ;
wire _07527_ ;
wire _07528_ ;
wire _07529_ ;
wire _07530_ ;
wire _07531_ ;
wire _07532_ ;
wire _07533_ ;
wire _07534_ ;
wire _07535_ ;
wire _07536_ ;
wire _07537_ ;
wire _07538_ ;
wire _07539_ ;
wire _07540_ ;
wire _07541_ ;
wire _07542_ ;
wire _07543_ ;
wire _07544_ ;
wire _07545_ ;
wire _07546_ ;
wire _07547_ ;
wire _07548_ ;
wire _07549_ ;
wire _07550_ ;
wire _07551_ ;
wire _07552_ ;
wire _07553_ ;
wire _07554_ ;
wire _07555_ ;
wire _07556_ ;
wire _07557_ ;
wire _07558_ ;
wire _07559_ ;
wire _07560_ ;
wire _07561_ ;
wire _07562_ ;
wire _07563_ ;
wire _07564_ ;
wire _07565_ ;
wire _07566_ ;
wire _07567_ ;
wire _07568_ ;
wire _07569_ ;
wire _07570_ ;
wire _07571_ ;
wire _07572_ ;
wire _07573_ ;
wire _07574_ ;
wire _07575_ ;
wire _07576_ ;
wire _07577_ ;
wire _07578_ ;
wire _07579_ ;
wire _07580_ ;
wire _07581_ ;
wire _07582_ ;
wire _07583_ ;
wire _07584_ ;
wire _07585_ ;
wire _07586_ ;
wire _07587_ ;
wire _07588_ ;
wire _07589_ ;
wire _07590_ ;
wire _07591_ ;
wire _07592_ ;
wire _07593_ ;
wire _07594_ ;
wire _07595_ ;
wire _07596_ ;
wire _07597_ ;
wire _07598_ ;
wire _07599_ ;
wire _07600_ ;
wire _07601_ ;
wire _07602_ ;
wire _07603_ ;
wire _07604_ ;
wire _07605_ ;
wire _07606_ ;
wire _07607_ ;
wire _07608_ ;
wire _07609_ ;
wire _07610_ ;
wire _07611_ ;
wire _07612_ ;
wire _07613_ ;
wire _07614_ ;
wire _07615_ ;
wire _07616_ ;
wire _07617_ ;
wire _07618_ ;
wire _07619_ ;
wire _07620_ ;
wire _07621_ ;
wire _07622_ ;
wire _07623_ ;
wire _07624_ ;
wire _07625_ ;
wire _07626_ ;
wire _07627_ ;
wire _07628_ ;
wire _07629_ ;
wire _07630_ ;
wire _07631_ ;
wire _07632_ ;
wire _07633_ ;
wire _07634_ ;
wire _07635_ ;
wire _07636_ ;
wire _07637_ ;
wire _07638_ ;
wire _07639_ ;
wire _07640_ ;
wire _07641_ ;
wire _07642_ ;
wire _07643_ ;
wire _07644_ ;
wire _07645_ ;
wire _07646_ ;
wire _07647_ ;
wire _07648_ ;
wire _07649_ ;
wire _07650_ ;
wire _07651_ ;
wire _07652_ ;
wire _07653_ ;
wire _07654_ ;
wire _07655_ ;
wire _07656_ ;
wire _07657_ ;
wire _07658_ ;
wire _07659_ ;
wire _07660_ ;
wire _07661_ ;
wire _07662_ ;
wire _07663_ ;
wire _07664_ ;
wire _07665_ ;
wire _07666_ ;
wire _07667_ ;
wire _07668_ ;
wire _07669_ ;
wire _07670_ ;
wire _07671_ ;
wire _07672_ ;
wire _07673_ ;
wire _07674_ ;
wire _07675_ ;
wire _07676_ ;
wire _07677_ ;
wire _07678_ ;
wire _07679_ ;
wire _07680_ ;
wire _07681_ ;
wire _07682_ ;
wire _07683_ ;
wire _07684_ ;
wire _07685_ ;
wire _07686_ ;
wire _07687_ ;
wire _07688_ ;
wire _07689_ ;
wire _07690_ ;
wire _07691_ ;
wire _07692_ ;
wire _07693_ ;
wire _07694_ ;
wire _07695_ ;
wire _07696_ ;
wire _07697_ ;
wire _07698_ ;
wire _07699_ ;
wire _07700_ ;
wire _07701_ ;
wire _07702_ ;
wire _07703_ ;
wire _07704_ ;
wire _07705_ ;
wire _07706_ ;
wire _07707_ ;
wire _07708_ ;
wire _07709_ ;
wire _07710_ ;
wire _07711_ ;
wire _07712_ ;
wire _07713_ ;
wire _07714_ ;
wire _07715_ ;
wire _07716_ ;
wire _07717_ ;
wire _07718_ ;
wire _07719_ ;
wire _07720_ ;
wire _07721_ ;
wire _07722_ ;
wire _07723_ ;
wire _07724_ ;
wire _07725_ ;
wire _07726_ ;
wire _07727_ ;
wire _07728_ ;
wire _07729_ ;
wire _07730_ ;
wire _07731_ ;
wire _07732_ ;
wire _07733_ ;
wire _07734_ ;
wire _07735_ ;
wire _07736_ ;
wire _07737_ ;
wire _07738_ ;
wire _07739_ ;
wire _07740_ ;
wire _07741_ ;
wire _07742_ ;
wire _07743_ ;
wire _07744_ ;
wire _07745_ ;
wire _07746_ ;
wire _07747_ ;
wire _07748_ ;
wire _07749_ ;
wire _07750_ ;
wire _07751_ ;
wire _07752_ ;
wire _07753_ ;
wire _07754_ ;
wire _07755_ ;
wire _07756_ ;
wire _07757_ ;
wire _07758_ ;
wire _07759_ ;
wire _07760_ ;
wire _07761_ ;
wire _07762_ ;
wire _07763_ ;
wire _07764_ ;
wire _07765_ ;
wire _07766_ ;
wire _07767_ ;
wire _07768_ ;
wire _07769_ ;
wire _07770_ ;
wire _07771_ ;
wire _07772_ ;
wire _07773_ ;
wire _07774_ ;
wire _07775_ ;
wire _07776_ ;
wire _07777_ ;
wire _07778_ ;
wire _07779_ ;
wire _07780_ ;
wire _07781_ ;
wire _07782_ ;
wire _07783_ ;
wire _07784_ ;
wire _07785_ ;
wire _07786_ ;
wire _07787_ ;
wire _07788_ ;
wire _07789_ ;
wire _07790_ ;
wire _07791_ ;
wire _07792_ ;
wire _07793_ ;
wire _07794_ ;
wire _07795_ ;
wire _07796_ ;
wire _07797_ ;
wire _07798_ ;
wire _07799_ ;
wire _07800_ ;
wire _07801_ ;
wire _07802_ ;
wire _07803_ ;
wire _07804_ ;
wire _07805_ ;
wire _07806_ ;
wire _07807_ ;
wire _07808_ ;
wire _07809_ ;
wire _07810_ ;
wire _07811_ ;
wire _07812_ ;
wire _07813_ ;
wire _07814_ ;
wire _07815_ ;
wire _07816_ ;
wire _07817_ ;
wire _07818_ ;
wire _07819_ ;
wire _07820_ ;
wire _07821_ ;
wire _07822_ ;
wire _07823_ ;
wire _07824_ ;
wire _07825_ ;
wire _07826_ ;
wire _07827_ ;
wire _07828_ ;
wire _07829_ ;
wire _07830_ ;
wire _07831_ ;
wire _07832_ ;
wire _07833_ ;
wire _07834_ ;
wire _07835_ ;
wire _07836_ ;
wire _07837_ ;
wire _07838_ ;
wire _07839_ ;
wire _07840_ ;
wire _07841_ ;
wire _07842_ ;
wire _07843_ ;
wire _07844_ ;
wire _07845_ ;
wire _07846_ ;
wire _07847_ ;
wire _07848_ ;
wire _07849_ ;
wire _07850_ ;
wire _07851_ ;
wire _07852_ ;
wire _07853_ ;
wire _07854_ ;
wire _07855_ ;
wire _07856_ ;
wire _07857_ ;
wire _07858_ ;
wire _07859_ ;
wire _07860_ ;
wire _07861_ ;
wire _07862_ ;
wire _07863_ ;
wire _07864_ ;
wire _07865_ ;
wire _07866_ ;
wire _07867_ ;
wire _07868_ ;
wire _07869_ ;
wire _07870_ ;
wire _07871_ ;
wire _07872_ ;
wire _07873_ ;
wire _07874_ ;
wire _07875_ ;
wire _07876_ ;
wire _07877_ ;
wire _07878_ ;
wire _07879_ ;
wire _07880_ ;
wire _07881_ ;
wire _07882_ ;
wire _07883_ ;
wire _07884_ ;
wire _07885_ ;
wire _07886_ ;
wire _07887_ ;
wire _07888_ ;
wire _07889_ ;
wire _07890_ ;
wire _07891_ ;
wire _07892_ ;
wire _07893_ ;
wire _07894_ ;
wire _07895_ ;
wire _07896_ ;
wire _07897_ ;
wire _07898_ ;
wire _07899_ ;
wire _07900_ ;
wire _07901_ ;
wire _07902_ ;
wire _07903_ ;
wire _07904_ ;
wire _07905_ ;
wire _07906_ ;
wire _07907_ ;
wire _07908_ ;
wire _07909_ ;
wire _07910_ ;
wire _07911_ ;
wire _07912_ ;
wire _07913_ ;
wire _07914_ ;
wire _07915_ ;
wire _07916_ ;
wire _07917_ ;
wire _07918_ ;
wire _07919_ ;
wire _07920_ ;
wire _07921_ ;
wire _07922_ ;
wire _07923_ ;
wire _07924_ ;
wire _07925_ ;
wire _07926_ ;
wire _07927_ ;
wire _07928_ ;
wire _07929_ ;
wire _07930_ ;
wire _07931_ ;
wire _07932_ ;
wire _07933_ ;
wire _07934_ ;
wire _07935_ ;
wire _07936_ ;
wire _07937_ ;
wire _07938_ ;
wire _07939_ ;
wire _07940_ ;
wire _07941_ ;
wire _07942_ ;
wire _07943_ ;
wire _07944_ ;
wire _07945_ ;
wire _07946_ ;
wire _07947_ ;
wire _07948_ ;
wire _07949_ ;
wire _07950_ ;
wire _07951_ ;
wire _07952_ ;
wire _07953_ ;
wire _07954_ ;
wire _07955_ ;
wire _07956_ ;
wire _07957_ ;
wire _07958_ ;
wire _07959_ ;
wire _07960_ ;
wire _07961_ ;
wire _07962_ ;
wire _07963_ ;
wire _07964_ ;
wire _07965_ ;
wire _07966_ ;
wire _07967_ ;
wire _07968_ ;
wire _07969_ ;
wire _07970_ ;
wire _07971_ ;
wire _07972_ ;
wire _07973_ ;
wire _07974_ ;
wire _07975_ ;
wire _07976_ ;
wire _07977_ ;
wire _07978_ ;
wire _07979_ ;
wire _07980_ ;
wire _07981_ ;
wire _07982_ ;
wire _07983_ ;
wire _07984_ ;
wire _07985_ ;
wire _07986_ ;
wire _07987_ ;
wire _07988_ ;
wire _07989_ ;
wire _07990_ ;
wire _07991_ ;
wire _07992_ ;
wire _07993_ ;
wire _07994_ ;
wire _07995_ ;
wire _07996_ ;
wire _07997_ ;
wire _07998_ ;
wire _07999_ ;
wire _08000_ ;
wire _08001_ ;
wire _08002_ ;
wire _08003_ ;
wire _08004_ ;
wire _08005_ ;
wire _08006_ ;
wire _08007_ ;
wire _08008_ ;
wire _08009_ ;
wire _08010_ ;
wire _08011_ ;
wire _08012_ ;
wire _08013_ ;
wire _08014_ ;
wire _08015_ ;
wire _08016_ ;
wire _08017_ ;
wire _08018_ ;
wire _08019_ ;
wire _08020_ ;
wire _08021_ ;
wire _08022_ ;
wire _08023_ ;
wire _08024_ ;
wire _08025_ ;
wire _08026_ ;
wire _08027_ ;
wire _08028_ ;
wire _08029_ ;
wire _08030_ ;
wire _08031_ ;
wire _08032_ ;
wire _08033_ ;
wire _08034_ ;
wire _08035_ ;
wire _08036_ ;
wire _08037_ ;
wire _08038_ ;
wire _08039_ ;
wire _08040_ ;
wire _08041_ ;
wire _08042_ ;
wire _08043_ ;
wire _08044_ ;
wire _08045_ ;
wire _08046_ ;
wire _08047_ ;
wire _08048_ ;
wire _08049_ ;
wire _08050_ ;
wire _08051_ ;
wire _08052_ ;
wire _08053_ ;
wire _08054_ ;
wire _08055_ ;
wire _08056_ ;
wire _08057_ ;
wire _08058_ ;
wire _08059_ ;
wire _08060_ ;
wire _08061_ ;
wire _08062_ ;
wire _08063_ ;
wire _08064_ ;
wire _08065_ ;
wire _08066_ ;
wire _08067_ ;
wire _08068_ ;
wire _08069_ ;
wire _08070_ ;
wire _08071_ ;
wire _08072_ ;
wire _08073_ ;
wire _08074_ ;
wire _08075_ ;
wire _08076_ ;
wire _08077_ ;
wire _08078_ ;
wire _08079_ ;
wire _08080_ ;
wire _08081_ ;
wire _08082_ ;
wire _08083_ ;
wire _08084_ ;
wire _08085_ ;
wire _08086_ ;
wire _08087_ ;
wire _08088_ ;
wire _08089_ ;
wire _08090_ ;
wire _08091_ ;
wire _08092_ ;
wire _08093_ ;
wire _08094_ ;
wire _08095_ ;
wire _08096_ ;
wire _08097_ ;
wire _08098_ ;
wire _08099_ ;
wire _08100_ ;
wire _08101_ ;
wire _08102_ ;
wire _08103_ ;
wire _08104_ ;
wire _08105_ ;
wire _08106_ ;
wire _08107_ ;
wire _08108_ ;
wire _08109_ ;
wire _08110_ ;
wire _08111_ ;
wire _08112_ ;
wire _08113_ ;
wire _08114_ ;
wire _08115_ ;
wire _08116_ ;
wire _08117_ ;
wire _08118_ ;
wire _08119_ ;
wire _08120_ ;
wire _08121_ ;
wire _08122_ ;
wire _08123_ ;
wire _08124_ ;
wire _08125_ ;
wire _08126_ ;
wire _08127_ ;
wire _08128_ ;
wire _08129_ ;
wire _08130_ ;
wire _08131_ ;
wire _08132_ ;
wire _08133_ ;
wire _08134_ ;
wire _08135_ ;
wire _08136_ ;
wire _08137_ ;
wire _08138_ ;
wire _08139_ ;
wire _08140_ ;
wire _08141_ ;
wire _08142_ ;
wire _08143_ ;
wire _08144_ ;
wire _08145_ ;
wire _08146_ ;
wire _08147_ ;
wire _08148_ ;
wire _08149_ ;
wire _08150_ ;
wire _08151_ ;
wire _08152_ ;
wire _08153_ ;
wire _08154_ ;
wire _08155_ ;
wire _08156_ ;
wire _08157_ ;
wire _08158_ ;
wire _08159_ ;
wire _08160_ ;
wire _08161_ ;
wire _08162_ ;
wire _08163_ ;
wire _08164_ ;
wire _08165_ ;
wire _08166_ ;
wire _08167_ ;
wire _08168_ ;
wire _08169_ ;
wire _08170_ ;
wire _08171_ ;
wire _08172_ ;
wire _08173_ ;
wire _08174_ ;
wire _08175_ ;
wire _08176_ ;
wire _08177_ ;
wire _08178_ ;
wire _08179_ ;
wire _08180_ ;
wire _08181_ ;
wire _08182_ ;
wire _08183_ ;
wire _08184_ ;
wire _08185_ ;
wire _08186_ ;
wire _08187_ ;
wire _08188_ ;
wire _08189_ ;
wire _08190_ ;
wire _08191_ ;
wire _08192_ ;
wire _08193_ ;
wire _08194_ ;
wire _08195_ ;
wire _08196_ ;
wire _08197_ ;
wire _08198_ ;
wire _08199_ ;
wire _08200_ ;
wire _08201_ ;
wire _08202_ ;
wire _08203_ ;
wire _08204_ ;
wire _08205_ ;
wire _08206_ ;
wire _08207_ ;
wire _08208_ ;
wire _08209_ ;
wire _08210_ ;
wire _08211_ ;
wire _08212_ ;
wire _08213_ ;
wire _08214_ ;
wire _08215_ ;
wire _08216_ ;
wire _08217_ ;
wire _08218_ ;
wire _08219_ ;
wire _08220_ ;
wire _08221_ ;
wire _08222_ ;
wire _08223_ ;
wire _08224_ ;
wire _08225_ ;
wire _08226_ ;
wire _08227_ ;
wire _08228_ ;
wire _08229_ ;
wire _08230_ ;
wire _08231_ ;
wire _08232_ ;
wire _08233_ ;
wire _08234_ ;
wire _08235_ ;
wire _08236_ ;
wire _08237_ ;
wire _08238_ ;
wire _08239_ ;
wire _08240_ ;
wire _08241_ ;
wire _08242_ ;
wire _08243_ ;
wire _08244_ ;
wire _08245_ ;
wire _08246_ ;
wire _08247_ ;
wire _08248_ ;
wire _08249_ ;
wire _08250_ ;
wire _08251_ ;
wire _08252_ ;
wire _08253_ ;
wire _08254_ ;
wire _08255_ ;
wire _08256_ ;
wire _08257_ ;
wire _08258_ ;
wire _08259_ ;
wire _08260_ ;
wire _08261_ ;
wire _08262_ ;
wire _08263_ ;
wire _08264_ ;
wire _08265_ ;
wire _08266_ ;
wire _08267_ ;
wire _08268_ ;
wire _08269_ ;
wire _08270_ ;
wire _08271_ ;
wire _08272_ ;
wire _08273_ ;
wire _08274_ ;
wire _08275_ ;
wire _08276_ ;
wire _08277_ ;
wire _08278_ ;
wire _08279_ ;
wire _08280_ ;
wire _08281_ ;
wire _08282_ ;
wire _08283_ ;
wire _08284_ ;
wire _08285_ ;
wire _08286_ ;
wire _08287_ ;
wire _08288_ ;
wire _08289_ ;
wire _08290_ ;
wire _08291_ ;
wire _08292_ ;
wire _08293_ ;
wire _08294_ ;
wire _08295_ ;
wire _08296_ ;
wire _08297_ ;
wire _08298_ ;
wire _08299_ ;
wire _08300_ ;
wire _08301_ ;
wire _08302_ ;
wire _08303_ ;
wire _08304_ ;
wire _08305_ ;
wire _08306_ ;
wire _08307_ ;
wire _08308_ ;
wire _08309_ ;
wire _08310_ ;
wire _08311_ ;
wire _08312_ ;
wire _08313_ ;
wire _08314_ ;
wire _08315_ ;
wire _08316_ ;
wire _08317_ ;
wire _08318_ ;
wire _08319_ ;
wire _08320_ ;
wire _08321_ ;
wire _08322_ ;
wire _08323_ ;
wire _08324_ ;
wire _08325_ ;
wire _08326_ ;
wire _08327_ ;
wire _08328_ ;
wire _08329_ ;
wire _08330_ ;
wire _08331_ ;
wire _08332_ ;
wire _08333_ ;
wire _08334_ ;
wire _08335_ ;
wire _08336_ ;
wire _08337_ ;
wire _08338_ ;
wire _08339_ ;
wire _08340_ ;
wire _08341_ ;
wire _08342_ ;
wire _08343_ ;
wire _08344_ ;
wire _08345_ ;
wire _08346_ ;
wire _08347_ ;
wire _08348_ ;
wire _08349_ ;
wire _08350_ ;
wire _08351_ ;
wire _08352_ ;
wire _08353_ ;
wire _08354_ ;
wire _08355_ ;
wire _08356_ ;
wire _08357_ ;
wire _08358_ ;
wire _08359_ ;
wire _08360_ ;
wire _08361_ ;
wire _08362_ ;
wire _08363_ ;
wire _08364_ ;
wire _08365_ ;
wire _08366_ ;
wire _08367_ ;
wire _08368_ ;
wire _08369_ ;
wire _08370_ ;
wire _08371_ ;
wire _08372_ ;
wire _08373_ ;
wire _08374_ ;
wire _08375_ ;
wire _08376_ ;
wire _08377_ ;
wire _08378_ ;
wire _08379_ ;
wire _08380_ ;
wire _08381_ ;
wire _08382_ ;
wire _08383_ ;
wire _08384_ ;
wire _08385_ ;
wire _08386_ ;
wire _08387_ ;
wire _08388_ ;
wire _08389_ ;
wire _08390_ ;
wire _08391_ ;
wire _08392_ ;
wire _08393_ ;
wire _08394_ ;
wire _08395_ ;
wire _08396_ ;
wire _08397_ ;
wire _08398_ ;
wire _08399_ ;
wire _08400_ ;
wire _08401_ ;
wire _08402_ ;
wire _08403_ ;
wire _08404_ ;
wire _08405_ ;
wire _08406_ ;
wire _08407_ ;
wire _08408_ ;
wire _08409_ ;
wire _08410_ ;
wire _08411_ ;
wire _08412_ ;
wire _08413_ ;
wire _08414_ ;
wire _08415_ ;
wire _08416_ ;
wire _08417_ ;
wire _08418_ ;
wire _08419_ ;
wire _08420_ ;
wire _08421_ ;
wire _08422_ ;
wire _08423_ ;
wire _08424_ ;
wire _08425_ ;
wire _08426_ ;
wire _08427_ ;
wire _08428_ ;
wire _08429_ ;
wire _08430_ ;
wire _08431_ ;
wire _08432_ ;
wire _08433_ ;
wire _08434_ ;
wire _08435_ ;
wire _08436_ ;
wire _08437_ ;
wire _08438_ ;
wire _08439_ ;
wire _08440_ ;
wire _08441_ ;
wire _08442_ ;
wire _08443_ ;
wire _08444_ ;
wire _08445_ ;
wire _08446_ ;
wire _08447_ ;
wire _08448_ ;
wire _08449_ ;
wire _08450_ ;
wire _08451_ ;
wire _08452_ ;
wire _08453_ ;
wire _08454_ ;
wire _08455_ ;
wire _08456_ ;
wire _08457_ ;
wire _08458_ ;
wire _08459_ ;
wire _08460_ ;
wire _08461_ ;
wire _08462_ ;
wire _08463_ ;
wire _08464_ ;
wire _08465_ ;
wire _08466_ ;
wire _08467_ ;
wire _08468_ ;
wire _08469_ ;
wire _08470_ ;
wire _08471_ ;
wire _08472_ ;
wire _08473_ ;
wire _08474_ ;
wire _08475_ ;
wire _08476_ ;
wire _08477_ ;
wire _08478_ ;
wire _08479_ ;
wire _08480_ ;
wire _08481_ ;
wire _08482_ ;
wire _08483_ ;
wire _08484_ ;
wire _08485_ ;
wire _08486_ ;
wire _08487_ ;
wire _08488_ ;
wire _08489_ ;
wire _08490_ ;
wire _08491_ ;
wire _08492_ ;
wire _08493_ ;
wire _08494_ ;
wire _08495_ ;
wire _08496_ ;
wire _08497_ ;
wire _08498_ ;
wire _08499_ ;
wire _08500_ ;
wire _08501_ ;
wire _08502_ ;
wire _08503_ ;
wire _08504_ ;
wire _08505_ ;
wire _08506_ ;
wire _08507_ ;
wire _08508_ ;
wire _08509_ ;
wire _08510_ ;
wire _08511_ ;
wire _08512_ ;
wire _08513_ ;
wire _08514_ ;
wire _08515_ ;
wire _08516_ ;
wire _08517_ ;
wire _08518_ ;
wire _08519_ ;
wire _08520_ ;
wire _08521_ ;
wire _08522_ ;
wire _08523_ ;
wire _08524_ ;
wire _08525_ ;
wire _08526_ ;
wire _08527_ ;
wire _08528_ ;
wire _08529_ ;
wire _08530_ ;
wire _08531_ ;
wire _08532_ ;
wire _08533_ ;
wire _08534_ ;
wire _08535_ ;
wire _08536_ ;
wire _08537_ ;
wire _08538_ ;
wire _08539_ ;
wire _08540_ ;
wire _08541_ ;
wire _08542_ ;
wire _08543_ ;
wire _08544_ ;
wire _08545_ ;
wire _08546_ ;
wire _08547_ ;
wire _08548_ ;
wire _08549_ ;
wire _08550_ ;
wire _08551_ ;
wire _08552_ ;
wire _08553_ ;
wire _08554_ ;
wire _08555_ ;
wire _08556_ ;
wire _08557_ ;
wire _08558_ ;
wire _08559_ ;
wire _08560_ ;
wire _08561_ ;
wire _08562_ ;
wire _08563_ ;
wire _08564_ ;
wire _08565_ ;
wire _08566_ ;
wire _08567_ ;
wire _08568_ ;
wire _08569_ ;
wire _08570_ ;
wire _08571_ ;
wire _08572_ ;
wire _08573_ ;
wire _08574_ ;
wire _08575_ ;
wire _08576_ ;
wire _08577_ ;
wire _08578_ ;
wire _08579_ ;
wire _08580_ ;
wire _08581_ ;
wire _08582_ ;
wire _08583_ ;
wire _08584_ ;
wire _08585_ ;
wire _08586_ ;
wire _08587_ ;
wire _08588_ ;
wire _08589_ ;
wire _08590_ ;
wire _08591_ ;
wire _08592_ ;
wire _08593_ ;
wire _08594_ ;
wire _08595_ ;
wire _08596_ ;
wire _08597_ ;
wire _08598_ ;
wire _08599_ ;
wire _08600_ ;
wire _08601_ ;
wire _08602_ ;
wire _08603_ ;
wire _08604_ ;
wire _08605_ ;
wire _08606_ ;
wire _08607_ ;
wire _08608_ ;
wire _08609_ ;
wire _08610_ ;
wire _08611_ ;
wire _08612_ ;
wire _08613_ ;
wire _08614_ ;
wire _08615_ ;
wire _08616_ ;
wire _08617_ ;
wire _08618_ ;
wire _08619_ ;
wire _08620_ ;
wire _08621_ ;
wire _08622_ ;
wire _08623_ ;
wire _08624_ ;
wire _08625_ ;
wire _08626_ ;
wire _08627_ ;
wire _08628_ ;
wire _08629_ ;
wire _08630_ ;
wire _08631_ ;
wire _08632_ ;
wire _08633_ ;
wire _08634_ ;
wire _08635_ ;
wire _08636_ ;
wire _08637_ ;
wire _08638_ ;
wire _08639_ ;
wire _08640_ ;
wire _08641_ ;
wire _08642_ ;
wire _08643_ ;
wire _08644_ ;
wire _08645_ ;
wire _08646_ ;
wire _08647_ ;
wire _08648_ ;
wire _08649_ ;
wire _08650_ ;
wire _08651_ ;
wire _08652_ ;
wire _08653_ ;
wire _08654_ ;
wire _08655_ ;
wire _08656_ ;
wire _08657_ ;
wire _08658_ ;
wire _08659_ ;
wire _08660_ ;
wire _08661_ ;
wire _08662_ ;
wire _08663_ ;
wire _08664_ ;
wire _08665_ ;
wire _08666_ ;
wire _08667_ ;
wire _08668_ ;
wire _08669_ ;
wire _08670_ ;
wire _08671_ ;
wire _08672_ ;
wire _08673_ ;
wire _08674_ ;
wire _08675_ ;
wire _08676_ ;
wire _08677_ ;
wire _08678_ ;
wire _08679_ ;
wire _08680_ ;
wire _08681_ ;
wire _08682_ ;
wire _08683_ ;
wire _08684_ ;
wire _08685_ ;
wire _08686_ ;
wire _08687_ ;
wire _08688_ ;
wire _08689_ ;
wire _08690_ ;
wire _08691_ ;
wire _08692_ ;
wire _08693_ ;
wire _08694_ ;
wire _08695_ ;
wire _08696_ ;
wire _08697_ ;
wire _08698_ ;
wire _08699_ ;
wire _08700_ ;
wire _08701_ ;
wire _08702_ ;
wire _08703_ ;
wire _08704_ ;
wire _08705_ ;
wire _08706_ ;
wire _08707_ ;
wire _08708_ ;
wire _08709_ ;
wire _08710_ ;
wire _08711_ ;
wire _08712_ ;
wire _08713_ ;
wire _08714_ ;
wire _08715_ ;
wire _08716_ ;
wire _08717_ ;
wire _08718_ ;
wire _08719_ ;
wire _08720_ ;
wire _08721_ ;
wire _08722_ ;
wire _08723_ ;
wire _08724_ ;
wire _08725_ ;
wire _08726_ ;
wire _08727_ ;
wire _08728_ ;
wire _08729_ ;
wire _08730_ ;
wire _08731_ ;
wire _08732_ ;
wire _08733_ ;
wire _08734_ ;
wire _08735_ ;
wire _08736_ ;
wire _08737_ ;
wire _08738_ ;
wire _08739_ ;
wire _08740_ ;
wire _08741_ ;
wire _08742_ ;
wire _08743_ ;
wire _08744_ ;
wire _08745_ ;
wire _08746_ ;
wire _08747_ ;
wire _08748_ ;
wire _08749_ ;
wire _08750_ ;
wire _08751_ ;
wire _08752_ ;
wire _08753_ ;
wire _08754_ ;
wire _08755_ ;
wire _08756_ ;
wire _08757_ ;
wire _08758_ ;
wire _08759_ ;
wire _08760_ ;
wire _08761_ ;
wire _08762_ ;
wire _08763_ ;
wire _08764_ ;
wire _08765_ ;
wire _08766_ ;
wire _08767_ ;
wire _08768_ ;
wire _08769_ ;
wire _08770_ ;
wire _08771_ ;
wire _08772_ ;
wire _08773_ ;
wire _08774_ ;
wire _08775_ ;
wire _08776_ ;
wire _08777_ ;
wire _08778_ ;
wire _08779_ ;
wire _08780_ ;
wire _08781_ ;
wire _08782_ ;
wire _08783_ ;
wire _08784_ ;
wire _08785_ ;
wire _08786_ ;
wire _08787_ ;
wire _08788_ ;
wire _08789_ ;
wire _08790_ ;
wire _08791_ ;
wire _08792_ ;
wire _08793_ ;
wire _08794_ ;
wire _08795_ ;
wire _08796_ ;
wire _08797_ ;
wire _08798_ ;
wire _08799_ ;
wire _08800_ ;
wire _08801_ ;
wire _08802_ ;
wire _08803_ ;
wire _08804_ ;
wire _08805_ ;
wire _08806_ ;
wire _08807_ ;
wire _08808_ ;
wire _08809_ ;
wire _08810_ ;
wire _08811_ ;
wire _08812_ ;
wire _08813_ ;
wire _08814_ ;
wire _08815_ ;
wire _08816_ ;
wire _08817_ ;
wire _08818_ ;
wire _08819_ ;
wire _08820_ ;
wire _08821_ ;
wire _08822_ ;
wire _08823_ ;
wire _08824_ ;
wire _08825_ ;
wire _08826_ ;
wire _08827_ ;
wire _08828_ ;
wire _08829_ ;
wire _08830_ ;
wire _08831_ ;
wire _08832_ ;
wire _08833_ ;
wire _08834_ ;
wire _08835_ ;
wire _08836_ ;
wire _08837_ ;
wire _08838_ ;
wire _08839_ ;
wire _08840_ ;
wire _08841_ ;
wire _08842_ ;
wire _08843_ ;
wire _08844_ ;
wire _08845_ ;
wire _08846_ ;
wire _08847_ ;
wire _08848_ ;
wire _08849_ ;
wire _08850_ ;
wire _08851_ ;
wire _08852_ ;
wire _08853_ ;
wire _08854_ ;
wire _08855_ ;
wire _08856_ ;
wire _08857_ ;
wire _08858_ ;
wire _08859_ ;
wire _08860_ ;
wire _08861_ ;
wire _08862_ ;
wire _08863_ ;
wire _08864_ ;
wire _08865_ ;
wire _08866_ ;
wire _08867_ ;
wire _08868_ ;
wire _08869_ ;
wire _08870_ ;
wire _08871_ ;
wire _08872_ ;
wire _08873_ ;
wire _08874_ ;
wire _08875_ ;
wire _08876_ ;
wire _08877_ ;
wire _08878_ ;
wire _08879_ ;
wire _08880_ ;
wire _08881_ ;
wire _08882_ ;
wire _08883_ ;
wire _08884_ ;
wire _08885_ ;
wire _08886_ ;
wire _08887_ ;
wire _08888_ ;
wire _08889_ ;
wire _08890_ ;
wire _08891_ ;
wire _08892_ ;
wire _08893_ ;
wire _08894_ ;
wire _08895_ ;
wire _08896_ ;
wire _08897_ ;
wire _08898_ ;
wire _08899_ ;
wire _08900_ ;
wire _08901_ ;
wire _08902_ ;
wire _08903_ ;
wire _08904_ ;
wire _08905_ ;
wire _08906_ ;
wire _08907_ ;
wire _08908_ ;
wire _08909_ ;
wire _08910_ ;
wire _08911_ ;
wire _08912_ ;
wire _08913_ ;
wire _08914_ ;
wire _08915_ ;
wire _08916_ ;
wire _08917_ ;
wire _08918_ ;
wire _08919_ ;
wire _08920_ ;
wire _08921_ ;
wire _08922_ ;
wire _08923_ ;
wire _08924_ ;
wire _08925_ ;
wire _08926_ ;
wire _08927_ ;
wire _08928_ ;
wire _08929_ ;
wire _08930_ ;
wire _08931_ ;
wire _08932_ ;
wire _08933_ ;
wire _08934_ ;
wire _08935_ ;
wire _08936_ ;
wire _08937_ ;
wire _08938_ ;
wire _08939_ ;
wire _08940_ ;
wire _08941_ ;
wire _08942_ ;
wire _08943_ ;
wire _08944_ ;
wire _08945_ ;
wire _08946_ ;
wire _08947_ ;
wire _08948_ ;
wire _08949_ ;
wire _08950_ ;
wire _08951_ ;
wire _08952_ ;
wire _08953_ ;
wire _08954_ ;
wire _08955_ ;
wire _08956_ ;
wire _08957_ ;
wire _08958_ ;
wire _08959_ ;
wire _08960_ ;
wire _08961_ ;
wire _08962_ ;
wire _08963_ ;
wire _08964_ ;
wire _08965_ ;
wire _08966_ ;
wire _08967_ ;
wire _08968_ ;
wire _08969_ ;
wire _08970_ ;
wire _08971_ ;
wire _08972_ ;
wire _08973_ ;
wire _08974_ ;
wire _08975_ ;
wire _08976_ ;
wire _08977_ ;
wire _08978_ ;
wire _08979_ ;
wire _08980_ ;
wire _08981_ ;
wire _08982_ ;
wire _08983_ ;
wire _08984_ ;
wire _08985_ ;
wire _08986_ ;
wire _08987_ ;
wire _08988_ ;
wire _08989_ ;
wire _08990_ ;
wire _08991_ ;
wire _08992_ ;
wire _08993_ ;
wire _08994_ ;
wire _08995_ ;
wire _08996_ ;
wire _08997_ ;
wire _08998_ ;
wire _08999_ ;
wire _09000_ ;
wire _09001_ ;
wire _09002_ ;
wire _09003_ ;
wire _09004_ ;
wire _09005_ ;
wire _09006_ ;
wire _09007_ ;
wire _09008_ ;
wire _09009_ ;
wire _09010_ ;
wire _09011_ ;
wire _09012_ ;
wire _09013_ ;
wire _09014_ ;
wire _09015_ ;
wire _09016_ ;
wire _09017_ ;
wire _09018_ ;
wire _09019_ ;
wire _09020_ ;
wire _09021_ ;
wire _09022_ ;
wire _09023_ ;
wire _09024_ ;
wire _09025_ ;
wire _09026_ ;
wire _09027_ ;
wire _09028_ ;
wire _09029_ ;
wire _09030_ ;
wire _09031_ ;
wire _09032_ ;
wire _09033_ ;
wire _09034_ ;
wire _09035_ ;
wire _09036_ ;
wire _09037_ ;
wire _09038_ ;
wire _09039_ ;
wire _09040_ ;
wire _09041_ ;
wire _09042_ ;
wire _09043_ ;
wire _09044_ ;
wire _09045_ ;
wire _09046_ ;
wire _09047_ ;
wire _09048_ ;
wire _09049_ ;
wire _09050_ ;
wire _09051_ ;
wire _09052_ ;
wire _09053_ ;
wire _09054_ ;
wire _09055_ ;
wire _09056_ ;
wire _09057_ ;
wire _09058_ ;
wire _09059_ ;
wire _09060_ ;
wire _09061_ ;
wire _09062_ ;
wire _09063_ ;
wire _09064_ ;
wire _09065_ ;
wire _09066_ ;
wire _09067_ ;
wire _09068_ ;
wire _09069_ ;
wire _09070_ ;
wire _09071_ ;
wire _09072_ ;
wire _09073_ ;
wire _09074_ ;
wire _09075_ ;
wire _09076_ ;
wire _09077_ ;
wire _09078_ ;
wire _09079_ ;
wire _09080_ ;
wire _09081_ ;
wire _09082_ ;
wire _09083_ ;
wire _09084_ ;
wire _09085_ ;
wire _09086_ ;
wire _09087_ ;
wire _09088_ ;
wire _09089_ ;
wire _09090_ ;
wire _09091_ ;
wire _09092_ ;
wire _09093_ ;
wire _09094_ ;
wire _09095_ ;
wire _09096_ ;
wire _09097_ ;
wire _09098_ ;
wire _09099_ ;
wire _09100_ ;
wire _09101_ ;
wire _09102_ ;
wire _09103_ ;
wire _09104_ ;
wire _09105_ ;
wire _09106_ ;
wire _09107_ ;
wire _09108_ ;
wire _09109_ ;
wire _09110_ ;
wire _09111_ ;
wire _09112_ ;
wire _09113_ ;
wire _09114_ ;
wire _09115_ ;
wire _09116_ ;
wire _09117_ ;
wire _09118_ ;
wire _09119_ ;
wire _09120_ ;
wire _09121_ ;
wire _09122_ ;
wire _09123_ ;
wire _09124_ ;
wire _09125_ ;
wire _09126_ ;
wire _09127_ ;
wire _09128_ ;
wire _09129_ ;
wire _09130_ ;
wire _09131_ ;
wire _09132_ ;
wire _09133_ ;
wire _09134_ ;
wire _09135_ ;
wire _09136_ ;
wire _09137_ ;
wire _09138_ ;
wire _09139_ ;
wire _09140_ ;
wire _09141_ ;
wire _09142_ ;
wire _09143_ ;
wire _09144_ ;
wire _09145_ ;
wire _09146_ ;
wire _09147_ ;
wire _09148_ ;
wire _09149_ ;
wire _09150_ ;
wire _09151_ ;
wire _09152_ ;
wire _09153_ ;
wire _09154_ ;
wire _09155_ ;
wire _09156_ ;
wire _09157_ ;
wire _09158_ ;
wire _09159_ ;
wire _09160_ ;
wire _09161_ ;
wire _09162_ ;
wire _09163_ ;
wire _09164_ ;
wire _09165_ ;
wire _09166_ ;
wire _09167_ ;
wire _09168_ ;
wire _09169_ ;
wire _09170_ ;
wire _09171_ ;
wire _09172_ ;
wire _09173_ ;
wire _09174_ ;
wire _09175_ ;
wire _09176_ ;
wire _09177_ ;
wire _09178_ ;
wire _09179_ ;
wire _09180_ ;
wire _09181_ ;
wire _09182_ ;
wire _09183_ ;
wire _09184_ ;
wire _09185_ ;
wire _09186_ ;
wire _09187_ ;
wire _09188_ ;
wire _09189_ ;
wire _09190_ ;
wire _09191_ ;
wire _09192_ ;
wire _09193_ ;
wire _09194_ ;
wire _09195_ ;
wire _09196_ ;
wire _09197_ ;
wire _09198_ ;
wire _09199_ ;
wire _09200_ ;
wire _09201_ ;
wire _09202_ ;
wire _09203_ ;
wire _09204_ ;
wire _09205_ ;
wire _09206_ ;
wire _09207_ ;
wire _09208_ ;
wire _09209_ ;
wire _09210_ ;
wire _09211_ ;
wire _09212_ ;
wire _09213_ ;
wire _09214_ ;
wire _09215_ ;
wire _09216_ ;
wire _09217_ ;
wire _09218_ ;
wire _09219_ ;
wire _09220_ ;
wire _09221_ ;
wire _09222_ ;
wire _09223_ ;
wire _09224_ ;
wire _09225_ ;
wire _09226_ ;
wire _09227_ ;
wire _09228_ ;
wire _09229_ ;
wire _09230_ ;
wire _09231_ ;
wire _09232_ ;
wire _09233_ ;
wire _09234_ ;
wire _09235_ ;
wire _09236_ ;
wire _09237_ ;
wire _09238_ ;
wire _09239_ ;
wire _09240_ ;
wire _09241_ ;
wire _09242_ ;
wire _09243_ ;
wire _09244_ ;
wire _09245_ ;
wire _09246_ ;
wire _09247_ ;
wire _09248_ ;
wire _09249_ ;
wire _09250_ ;
wire _09251_ ;
wire _09252_ ;
wire _09253_ ;
wire _09254_ ;
wire _09255_ ;
wire _09256_ ;
wire _09257_ ;
wire _09258_ ;
wire _09259_ ;
wire _09260_ ;
wire _09261_ ;
wire _09262_ ;
wire _09263_ ;
wire _09264_ ;
wire _09265_ ;
wire _09266_ ;
wire _09267_ ;
wire _09268_ ;
wire _09269_ ;
wire _09270_ ;
wire _09271_ ;
wire _09272_ ;
wire _09273_ ;
wire _09274_ ;
wire _09275_ ;
wire _09276_ ;
wire _09277_ ;
wire _09278_ ;
wire _09279_ ;
wire _09280_ ;
wire _09281_ ;
wire _09282_ ;
wire _09283_ ;
wire _09284_ ;
wire _09285_ ;
wire _09286_ ;
wire _09287_ ;
wire _09288_ ;
wire _09289_ ;
wire _09290_ ;
wire _09291_ ;
wire _09292_ ;
wire _09293_ ;
wire _09294_ ;
wire _09295_ ;
wire _09296_ ;
wire _09297_ ;
wire _09298_ ;
wire _09299_ ;
wire _09300_ ;
wire _09301_ ;
wire _09302_ ;
wire _09303_ ;
wire _09304_ ;
wire _09305_ ;
wire _09306_ ;
wire _09307_ ;
wire _09308_ ;
wire _09309_ ;
wire _09310_ ;
wire _09311_ ;
wire _09312_ ;
wire _09313_ ;
wire _09314_ ;
wire _09315_ ;
wire _09316_ ;
wire _09317_ ;
wire _09318_ ;
wire _09319_ ;
wire _09320_ ;
wire _09321_ ;
wire _09322_ ;
wire _09323_ ;
wire _09324_ ;
wire _09325_ ;
wire _09326_ ;
wire _09327_ ;
wire _09328_ ;
wire _09329_ ;
wire _09330_ ;
wire _09331_ ;
wire _09332_ ;
wire _09333_ ;
wire _09334_ ;
wire _09335_ ;
wire _09336_ ;
wire _09337_ ;
wire _09338_ ;
wire _09339_ ;
wire _09340_ ;
wire _09341_ ;
wire _09342_ ;
wire _09343_ ;
wire _09344_ ;
wire _09345_ ;
wire _09346_ ;
wire _09347_ ;
wire _09348_ ;
wire _09349_ ;
wire _09350_ ;
wire _09351_ ;
wire _09352_ ;
wire _09353_ ;
wire _09354_ ;
wire _09355_ ;
wire _09356_ ;
wire _09357_ ;
wire _09358_ ;
wire _09359_ ;
wire _09360_ ;
wire _09361_ ;
wire _09362_ ;
wire _09363_ ;
wire _09364_ ;
wire _09365_ ;
wire _09366_ ;
wire _09367_ ;
wire _09368_ ;
wire _09369_ ;
wire _09370_ ;
wire _09371_ ;
wire _09372_ ;
wire _09373_ ;
wire _09374_ ;
wire _09375_ ;
wire _09376_ ;
wire _09377_ ;
wire _09378_ ;
wire _09379_ ;
wire _09380_ ;
wire _09381_ ;
wire _09382_ ;
wire _09383_ ;
wire _09384_ ;
wire _09385_ ;
wire _09386_ ;
wire _09387_ ;
wire _09388_ ;
wire _09389_ ;
wire _09390_ ;
wire _09391_ ;
wire _09392_ ;
wire _09393_ ;
wire _09394_ ;
wire _09395_ ;
wire _09396_ ;
wire _09397_ ;
wire _09398_ ;
wire _09399_ ;
wire _09400_ ;
wire _09401_ ;
wire _09402_ ;
wire _09403_ ;
wire _09404_ ;
wire _09405_ ;
wire _09406_ ;
wire _09407_ ;
wire _09408_ ;
wire _09409_ ;
wire _09410_ ;
wire _09411_ ;
wire _09412_ ;
wire _09413_ ;
wire _09414_ ;
wire _09415_ ;
wire _09416_ ;
wire _09417_ ;
wire _09418_ ;
wire _09419_ ;
wire _09420_ ;
wire _09421_ ;
wire _09422_ ;
wire _09423_ ;
wire _09424_ ;
wire _09425_ ;
wire _09426_ ;
wire _09427_ ;
wire _09428_ ;
wire _09429_ ;
wire _09430_ ;
wire _09431_ ;
wire _09432_ ;
wire _09433_ ;
wire _09434_ ;
wire _09435_ ;
wire _09436_ ;
wire _09437_ ;
wire _09438_ ;
wire _09439_ ;
wire _09440_ ;
wire _09441_ ;
wire _09442_ ;
wire _09443_ ;
wire _09444_ ;
wire _09445_ ;
wire _09446_ ;
wire _09447_ ;
wire _09448_ ;
wire _09449_ ;
wire _09450_ ;
wire _09451_ ;
wire _09452_ ;
wire _09453_ ;
wire _09454_ ;
wire _09455_ ;
wire _09456_ ;
wire _09457_ ;
wire _09458_ ;
wire _09459_ ;
wire _09460_ ;
wire _09461_ ;
wire _09462_ ;
wire _09463_ ;
wire _09464_ ;
wire _09465_ ;
wire _09466_ ;
wire _09467_ ;
wire _09468_ ;
wire _09469_ ;
wire _09470_ ;
wire _09471_ ;
wire _09472_ ;
wire _09473_ ;
wire _09474_ ;
wire _09475_ ;
wire _09476_ ;
wire _09477_ ;
wire _09478_ ;
wire _09479_ ;
wire _09480_ ;
wire _09481_ ;
wire _09482_ ;
wire _09483_ ;
wire _09484_ ;
wire _09485_ ;
wire _09486_ ;
wire _09487_ ;
wire _09488_ ;
wire _09489_ ;
wire _09490_ ;
wire _09491_ ;
wire _09492_ ;
wire _09493_ ;
wire _09494_ ;
wire _09495_ ;
wire _09496_ ;
wire _09497_ ;
wire _09498_ ;
wire _09499_ ;
wire _09500_ ;
wire _09501_ ;
wire _09502_ ;
wire _09503_ ;
wire _09504_ ;
wire _09505_ ;
wire _09506_ ;
wire _09507_ ;
wire _09508_ ;
wire _09509_ ;
wire _09510_ ;
wire _09511_ ;
wire _09512_ ;
wire _09513_ ;
wire _09514_ ;
wire _09515_ ;
wire _09516_ ;
wire _09517_ ;
wire _09518_ ;
wire _09519_ ;
wire _09520_ ;
wire _09521_ ;
wire _09522_ ;
wire _09523_ ;
wire _09524_ ;
wire _09525_ ;
wire _09526_ ;
wire _09527_ ;
wire _09528_ ;
wire _09529_ ;
wire _09530_ ;
wire _09531_ ;
wire _09532_ ;
wire _09533_ ;
wire _09534_ ;
wire _09535_ ;
wire _09536_ ;
wire _09537_ ;
wire _09538_ ;
wire _09539_ ;
wire _09540_ ;
wire _09541_ ;
wire _09542_ ;
wire _09543_ ;
wire _09544_ ;
wire _09545_ ;
wire _09546_ ;
wire _09547_ ;
wire _09548_ ;
wire _09549_ ;
wire _09550_ ;
wire _09551_ ;
wire _09552_ ;
wire _09553_ ;
wire _09554_ ;
wire _09555_ ;
wire _09556_ ;
wire _09557_ ;
wire _09558_ ;
wire _09559_ ;
wire _09560_ ;
wire _09561_ ;
wire _09562_ ;
wire _09563_ ;
wire _09564_ ;
wire _09565_ ;
wire _09566_ ;
wire _09567_ ;
wire _09568_ ;
wire _09569_ ;
wire _09570_ ;
wire _09571_ ;
wire _09572_ ;
wire _09573_ ;
wire _09574_ ;
wire _09575_ ;
wire _09576_ ;
wire _09577_ ;
wire _09578_ ;
wire _09579_ ;
wire _09580_ ;
wire _09581_ ;
wire _09582_ ;
wire _09583_ ;
wire _09584_ ;
wire _09585_ ;
wire _09586_ ;
wire _09587_ ;
wire _09588_ ;
wire _09589_ ;
wire _09590_ ;
wire _09591_ ;
wire _09592_ ;
wire _09593_ ;
wire _09594_ ;
wire _09595_ ;
wire _09596_ ;
wire _09597_ ;
wire _09598_ ;
wire _09599_ ;
wire _09600_ ;
wire _09601_ ;
wire _09602_ ;
wire _09603_ ;
wire _09604_ ;
wire _09605_ ;
wire _09606_ ;
wire _09607_ ;
wire _09608_ ;
wire _09609_ ;
wire _09610_ ;
wire _09611_ ;
wire _09612_ ;
wire _09613_ ;
wire _09614_ ;
wire _09615_ ;
wire _09616_ ;
wire _09617_ ;
wire _09618_ ;
wire _09619_ ;
wire _09620_ ;
wire _09621_ ;
wire _09622_ ;
wire _09623_ ;
wire _09624_ ;
wire _09625_ ;
wire _09626_ ;
wire _09627_ ;
wire _09628_ ;
wire _09629_ ;
wire _09630_ ;
wire _09631_ ;
wire _09632_ ;
wire _09633_ ;
wire _09634_ ;
wire _09635_ ;
wire _09636_ ;
wire _09637_ ;
wire _09638_ ;
wire _09639_ ;
wire _09640_ ;
wire _09641_ ;
wire _09642_ ;
wire _09643_ ;
wire _09644_ ;
wire _09645_ ;
wire _09646_ ;
wire _09647_ ;
wire _09648_ ;
wire _09649_ ;
wire _09650_ ;
wire _09651_ ;
wire _09652_ ;
wire _09653_ ;
wire _09654_ ;
wire _09655_ ;
wire _09656_ ;
wire _09657_ ;
wire _09658_ ;
wire _09659_ ;
wire _09660_ ;
wire _09661_ ;
wire _09662_ ;
wire _09663_ ;
wire _09664_ ;
wire _09665_ ;
wire _09666_ ;
wire _09667_ ;
wire _09668_ ;
wire _09669_ ;
wire _09670_ ;
wire _09671_ ;
wire _09672_ ;
wire _09673_ ;
wire _09674_ ;
wire _09675_ ;
wire _09676_ ;
wire _09677_ ;
wire _09678_ ;
wire _09679_ ;
wire _09680_ ;
wire _09681_ ;
wire _09682_ ;
wire _09683_ ;
wire _09684_ ;
wire _09685_ ;
wire _09686_ ;
wire _09687_ ;
wire _09688_ ;
wire _09689_ ;
wire _09690_ ;
wire _09691_ ;
wire _09692_ ;
wire _09693_ ;
wire _09694_ ;
wire _09695_ ;
wire _09696_ ;
wire _09697_ ;
wire _09698_ ;
wire _09699_ ;
wire _09700_ ;
wire _09701_ ;
wire _09702_ ;
wire _09703_ ;
wire _09704_ ;
wire _09705_ ;
wire _09706_ ;
wire _09707_ ;
wire _09708_ ;
wire _09709_ ;
wire _09710_ ;
wire _09711_ ;
wire _09712_ ;
wire _09713_ ;
wire _09714_ ;
wire _09715_ ;
wire _09716_ ;
wire _09717_ ;
wire _09718_ ;
wire _09719_ ;
wire _09720_ ;
wire _09721_ ;
wire _09722_ ;
wire _09723_ ;
wire _09724_ ;
wire _09725_ ;
wire _09726_ ;
wire _09727_ ;
wire _09728_ ;
wire _09729_ ;
wire _09730_ ;
wire _09731_ ;
wire _09732_ ;
wire _09733_ ;
wire _09734_ ;
wire _09735_ ;
wire _09736_ ;
wire _09737_ ;
wire _09738_ ;
wire _09739_ ;
wire _09740_ ;
wire _09741_ ;
wire _09742_ ;
wire _09743_ ;
wire _09744_ ;
wire _09745_ ;
wire _09746_ ;
wire _09747_ ;
wire _09748_ ;
wire _09749_ ;
wire _09750_ ;
wire _09751_ ;
wire _09752_ ;
wire _09753_ ;
wire _09754_ ;
wire _09755_ ;
wire _09756_ ;
wire _09757_ ;
wire _09758_ ;
wire _09759_ ;
wire _09760_ ;
wire _09761_ ;
wire _09762_ ;
wire _09763_ ;
wire _09764_ ;
wire _09765_ ;
wire _09766_ ;
wire _09767_ ;
wire _09768_ ;
wire _09769_ ;
wire _09770_ ;
wire _09771_ ;
wire _09772_ ;
wire _09773_ ;
wire _09774_ ;
wire _09775_ ;
wire _09776_ ;
wire _09777_ ;
wire _09778_ ;
wire _09779_ ;
wire _09780_ ;
wire _09781_ ;
wire _09782_ ;
wire _09783_ ;
wire _09784_ ;
wire _09785_ ;
wire _09786_ ;
wire _09787_ ;
wire _09788_ ;
wire _09789_ ;
wire _09790_ ;
wire _09791_ ;
wire _09792_ ;
wire _09793_ ;
wire _09794_ ;
wire _09795_ ;
wire _09796_ ;
wire _09797_ ;
wire _09798_ ;
wire _09799_ ;
wire _09800_ ;
wire _09801_ ;
wire _09802_ ;
wire _09803_ ;
wire _09804_ ;
wire _09805_ ;
wire _09806_ ;
wire _09807_ ;
wire _09808_ ;
wire _09809_ ;
wire _09810_ ;
wire _09811_ ;
wire _09812_ ;
wire _09813_ ;
wire _09814_ ;
wire _09815_ ;
wire _09816_ ;
wire _09817_ ;
wire _09818_ ;
wire _09819_ ;
wire _09820_ ;
wire _09821_ ;
wire _09822_ ;
wire _09823_ ;
wire _09824_ ;
wire _09825_ ;
wire _09826_ ;
wire _09827_ ;
wire _09828_ ;
wire _09829_ ;
wire _09830_ ;
wire _09831_ ;
wire _09832_ ;
wire _09833_ ;
wire _09834_ ;
wire _09835_ ;
wire _09836_ ;
wire _09837_ ;
wire _09838_ ;
wire _09839_ ;
wire _09840_ ;
wire _09841_ ;
wire _09842_ ;
wire _09843_ ;
wire _09844_ ;
wire _09845_ ;
wire _09846_ ;
wire _09847_ ;
wire _09848_ ;
wire _09849_ ;
wire _09850_ ;
wire _09851_ ;
wire _09852_ ;
wire _09853_ ;
wire _09854_ ;
wire _09855_ ;
wire _09856_ ;
wire _09857_ ;
wire _09858_ ;
wire _09859_ ;
wire _09860_ ;
wire _09861_ ;
wire _09862_ ;
wire _09863_ ;
wire _09864_ ;
wire _09865_ ;
wire _09866_ ;
wire _09867_ ;
wire _09868_ ;
wire _09869_ ;
wire _09870_ ;
wire _09871_ ;
wire _09872_ ;
wire _09873_ ;
wire _09874_ ;
wire _09875_ ;
wire _09876_ ;
wire _09877_ ;
wire _09878_ ;
wire _09879_ ;
wire _09880_ ;
wire _09881_ ;
wire _09882_ ;
wire _09883_ ;
wire _09884_ ;
wire _09885_ ;
wire _09886_ ;
wire _09887_ ;
wire _09888_ ;
wire _09889_ ;
wire _09890_ ;
wire _09891_ ;
wire _09892_ ;
wire _09893_ ;
wire _09894_ ;
wire _09895_ ;
wire _09896_ ;
wire _09897_ ;
wire _09898_ ;
wire _09899_ ;
wire _09900_ ;
wire _09901_ ;
wire _09902_ ;
wire _09903_ ;
wire _09904_ ;
wire _09905_ ;
wire _09906_ ;
wire _09907_ ;
wire _09908_ ;
wire _09909_ ;
wire _09910_ ;
wire _09911_ ;
wire _09912_ ;
wire _09913_ ;
wire _09914_ ;
wire _09915_ ;
wire _09916_ ;
wire _09917_ ;
wire _09918_ ;
wire _09919_ ;
wire _09920_ ;
wire _09921_ ;
wire _09922_ ;
wire _09923_ ;
wire _09924_ ;
wire _09925_ ;
wire _09926_ ;
wire _09927_ ;
wire _09928_ ;
wire _09929_ ;
wire _09930_ ;
wire _09931_ ;
wire _09932_ ;
wire _09933_ ;
wire _09934_ ;
wire _09935_ ;
wire _09936_ ;
wire _09937_ ;
wire _09938_ ;
wire _09939_ ;
wire _09940_ ;
wire _09941_ ;
wire _09942_ ;
wire _09943_ ;
wire _09944_ ;
wire _09945_ ;
wire _09946_ ;
wire _09947_ ;
wire _09948_ ;
wire _09949_ ;
wire _09950_ ;
wire _09951_ ;
wire _09952_ ;
wire _09953_ ;
wire _09954_ ;
wire _09955_ ;
wire _09956_ ;
wire _09957_ ;
wire _09958_ ;
wire _09959_ ;
wire _09960_ ;
wire _09961_ ;
wire _09962_ ;
wire _09963_ ;
wire _09964_ ;
wire _09965_ ;
wire _09966_ ;
wire _09967_ ;
wire _09968_ ;
wire _09969_ ;
wire _09970_ ;
wire _09971_ ;
wire _09972_ ;
wire _09973_ ;
wire _09974_ ;
wire _09975_ ;
wire _09976_ ;
wire _09977_ ;
wire _09978_ ;
wire _09979_ ;
wire _09980_ ;
wire _09981_ ;
wire _09982_ ;
wire _09983_ ;
wire _09984_ ;
wire _09985_ ;
wire _09986_ ;
wire _09987_ ;
wire _09988_ ;
wire _09989_ ;
wire _09990_ ;
wire _09991_ ;
wire _09992_ ;
wire _09993_ ;
wire _09994_ ;
wire _09995_ ;
wire _09996_ ;
wire _09997_ ;
wire _09998_ ;
wire _09999_ ;
wire _10000_ ;
wire _10001_ ;
wire _10002_ ;
wire _10003_ ;
wire _10004_ ;
wire _10005_ ;
wire _10006_ ;
wire _10007_ ;
wire _10008_ ;
wire _10009_ ;
wire _10010_ ;
wire _10011_ ;
wire _10012_ ;
wire _10013_ ;
wire _10014_ ;
wire _10015_ ;
wire _10016_ ;
wire _10017_ ;
wire _10018_ ;
wire _10019_ ;
wire _10020_ ;
wire _10021_ ;
wire _10022_ ;
wire _10023_ ;
wire _10024_ ;
wire _10025_ ;
wire _10026_ ;
wire _10027_ ;
wire _10028_ ;
wire _10029_ ;
wire _10030_ ;
wire _10031_ ;
wire _10032_ ;
wire _10033_ ;
wire _10034_ ;
wire _10035_ ;
wire _10036_ ;
wire _10037_ ;
wire _10038_ ;
wire _10039_ ;
wire _10040_ ;
wire _10041_ ;
wire _10042_ ;
wire _10043_ ;
wire _10044_ ;
wire _10045_ ;
wire _10046_ ;
wire _10047_ ;
wire _10048_ ;
wire _10049_ ;
wire _10050_ ;
wire _10051_ ;
wire _10052_ ;
wire _10053_ ;
wire _10054_ ;
wire _10055_ ;
wire _10056_ ;
wire _10057_ ;
wire _10058_ ;
wire _10059_ ;
wire _10060_ ;
wire _10061_ ;
wire _10062_ ;
wire _10063_ ;
wire _10064_ ;
wire _10065_ ;
wire _10066_ ;
wire _10067_ ;
wire _10068_ ;
wire _10069_ ;
wire _10070_ ;
wire _10071_ ;
wire _10072_ ;
wire _10073_ ;
wire _10074_ ;
wire _10075_ ;
wire _10076_ ;
wire _10077_ ;
wire _10078_ ;
wire _10079_ ;
wire _10080_ ;
wire _10081_ ;
wire _10082_ ;
wire _10083_ ;
wire _10084_ ;
wire _10085_ ;
wire _10086_ ;
wire _10087_ ;
wire _10088_ ;
wire _10089_ ;
wire _10090_ ;
wire _10091_ ;
wire _10092_ ;
wire _10093_ ;
wire _10094_ ;
wire _10095_ ;
wire _10096_ ;
wire _10097_ ;
wire _10098_ ;
wire _10099_ ;
wire _10100_ ;
wire _10101_ ;
wire _10102_ ;
wire _10103_ ;
wire _10104_ ;
wire _10105_ ;
wire _10106_ ;
wire _10107_ ;
wire _10108_ ;
wire _10109_ ;
wire _10110_ ;
wire _10111_ ;
wire _10112_ ;
wire _10113_ ;
wire _10114_ ;
wire _10115_ ;
wire _10116_ ;
wire _10117_ ;
wire _10118_ ;
wire _10119_ ;
wire _10120_ ;
wire _10121_ ;
wire _10122_ ;
wire _10123_ ;
wire _10124_ ;
wire _10125_ ;
wire _10126_ ;
wire _10127_ ;
wire _10128_ ;
wire _10129_ ;
wire _10130_ ;
wire _10131_ ;
wire _10132_ ;
wire _10133_ ;
wire _10134_ ;
wire _10135_ ;
wire _10136_ ;
wire _10137_ ;
wire _10138_ ;
wire _10139_ ;
wire _10140_ ;
wire _10141_ ;
wire _10142_ ;
wire _10143_ ;
wire _10144_ ;
wire _10145_ ;
wire _10146_ ;
wire _10147_ ;
wire _10148_ ;
wire _10149_ ;
wire _10150_ ;
wire _10151_ ;
wire _10152_ ;
wire _10153_ ;
wire _10154_ ;
wire _10155_ ;
wire _10156_ ;
wire _10157_ ;
wire _10158_ ;
wire _10159_ ;
wire _10160_ ;
wire _10161_ ;
wire _10162_ ;
wire _10163_ ;
wire _10164_ ;
wire _10165_ ;
wire _10166_ ;
wire _10167_ ;
wire _10168_ ;
wire _10169_ ;
wire _10170_ ;
wire _10171_ ;
wire _10172_ ;
wire _10173_ ;
wire _10174_ ;
wire _10175_ ;
wire _10176_ ;
wire _10177_ ;
wire _10178_ ;
wire _10179_ ;
wire _10180_ ;
wire _10181_ ;
wire _10182_ ;
wire _10183_ ;
wire _10184_ ;
wire _10185_ ;
wire _10186_ ;
wire _10187_ ;
wire _10188_ ;
wire _10189_ ;
wire _10190_ ;
wire _10191_ ;
wire _10192_ ;
wire _10193_ ;
wire _10194_ ;
wire _10195_ ;
wire _10196_ ;
wire _10197_ ;
wire _10198_ ;
wire _10199_ ;
wire _10200_ ;
wire _10201_ ;
wire _10202_ ;
wire _10203_ ;
wire _10204_ ;
wire _10205_ ;
wire _10206_ ;
wire _10207_ ;
wire _10208_ ;
wire _10209_ ;
wire _10210_ ;
wire _10211_ ;
wire _10212_ ;
wire _10213_ ;
wire _10214_ ;
wire _10215_ ;
wire _10216_ ;
wire _10217_ ;
wire _10218_ ;
wire _10219_ ;
wire _10220_ ;
wire _10221_ ;
wire _10222_ ;
wire _10223_ ;
wire _10224_ ;
wire _10225_ ;
wire _10226_ ;
wire _10227_ ;
wire _10228_ ;
wire _10229_ ;
wire _10230_ ;
wire _10231_ ;
wire _10232_ ;
wire _10233_ ;
wire _10234_ ;
wire _10235_ ;
wire _10236_ ;
wire _10237_ ;
wire _10238_ ;
wire _10239_ ;
wire _10240_ ;
wire _10241_ ;
wire _10242_ ;
wire _10243_ ;
wire _10244_ ;
wire _10245_ ;
wire _10246_ ;
wire _10247_ ;
wire _10248_ ;
wire _10249_ ;
wire _10250_ ;
wire _10251_ ;
wire _10252_ ;
wire _10253_ ;
wire _10254_ ;
wire _10255_ ;
wire _10256_ ;
wire _10257_ ;
wire _10258_ ;
wire _10259_ ;
wire _10260_ ;
wire _10261_ ;
wire _10262_ ;
wire _10263_ ;
wire _10264_ ;
wire _10265_ ;
wire _10266_ ;
wire _10267_ ;
wire _10268_ ;
wire _10269_ ;
wire _10270_ ;
wire _10271_ ;
wire _10272_ ;
wire _10273_ ;
wire _10274_ ;
wire _10275_ ;
wire _10276_ ;
wire _10277_ ;
wire _10278_ ;
wire _10279_ ;
wire _10280_ ;
wire _10281_ ;
wire _10282_ ;
wire _10283_ ;
wire _10284_ ;
wire _10285_ ;
wire _10286_ ;
wire _10287_ ;
wire _10288_ ;
wire _10289_ ;
wire _10290_ ;
wire _10291_ ;
wire _10292_ ;
wire _10293_ ;
wire _10294_ ;
wire _10295_ ;
wire _10296_ ;
wire _10297_ ;
wire _10298_ ;
wire _10299_ ;
wire _10300_ ;
wire _10301_ ;
wire _10302_ ;
wire _10303_ ;
wire _10304_ ;
wire _10305_ ;
wire _10306_ ;
wire _10307_ ;
wire _10308_ ;
wire _10309_ ;
wire _10310_ ;
wire _10311_ ;
wire _10312_ ;
wire _10313_ ;
wire _10314_ ;
wire _10315_ ;
wire _10316_ ;
wire _10317_ ;
wire _10318_ ;
wire _10319_ ;
wire _10320_ ;
wire _10321_ ;
wire _10322_ ;
wire _10323_ ;
wire _10324_ ;
wire _10325_ ;
wire _10326_ ;
wire _10327_ ;
wire _10328_ ;
wire _10329_ ;
wire _10330_ ;
wire _10331_ ;
wire _10332_ ;
wire _10333_ ;
wire _10334_ ;
wire _10335_ ;
wire _10336_ ;
wire _10337_ ;
wire _10338_ ;
wire _10339_ ;
wire _10340_ ;
wire _10341_ ;
wire _10342_ ;
wire _10343_ ;
wire _10344_ ;
wire _10345_ ;
wire _10346_ ;
wire _10347_ ;
wire _10348_ ;
wire _10349_ ;
wire _10350_ ;
wire _10351_ ;
wire _10352_ ;
wire _10353_ ;
wire _10354_ ;
wire _10355_ ;
wire _10356_ ;
wire _10357_ ;
wire _10358_ ;
wire _10359_ ;
wire _10360_ ;
wire _10361_ ;
wire _10362_ ;
wire _10363_ ;
wire _10364_ ;
wire _10365_ ;
wire _10366_ ;
wire _10367_ ;
wire _10368_ ;
wire _10369_ ;
wire _10370_ ;
wire _10371_ ;
wire _10372_ ;
wire _10373_ ;
wire _10374_ ;
wire _10375_ ;
wire _10376_ ;
wire _10377_ ;
wire _10378_ ;
wire _10379_ ;
wire _10380_ ;
wire _10381_ ;
wire _10382_ ;
wire _10383_ ;
wire _10384_ ;
wire _10385_ ;
wire _10386_ ;
wire _10387_ ;
wire _10388_ ;
wire _10389_ ;
wire _10390_ ;
wire _10391_ ;
wire _10392_ ;
wire _10393_ ;
wire _10394_ ;
wire _10395_ ;
wire _10396_ ;
wire _10397_ ;
wire _10398_ ;
wire _10399_ ;
wire _10400_ ;
wire _10401_ ;
wire _10402_ ;
wire _10403_ ;
wire _10404_ ;
wire _10405_ ;
wire _10406_ ;
wire _10407_ ;
wire _10408_ ;
wire _10409_ ;
wire _10410_ ;
wire _10411_ ;
wire _10412_ ;
wire _10413_ ;
wire _10414_ ;
wire _10415_ ;
wire _10416_ ;
wire _10417_ ;
wire _10418_ ;
wire _10419_ ;
wire _10420_ ;
wire _10421_ ;
wire _10422_ ;
wire _10423_ ;
wire _10424_ ;
wire _10425_ ;
wire _10426_ ;
wire _10427_ ;
wire _10428_ ;
wire _10429_ ;
wire _10430_ ;
wire _10431_ ;
wire _10432_ ;
wire _10433_ ;
wire _10434_ ;
wire _10435_ ;
wire _10436_ ;
wire _10437_ ;
wire _10438_ ;
wire _10439_ ;
wire _10440_ ;
wire _10441_ ;
wire _10442_ ;
wire _10443_ ;
wire _10444_ ;
wire _10445_ ;
wire _10446_ ;
wire _10447_ ;
wire _10448_ ;
wire _10449_ ;
wire _10450_ ;
wire _10451_ ;
wire _10452_ ;
wire _10453_ ;
wire _10454_ ;
wire _10455_ ;
wire _10456_ ;
wire _10457_ ;
wire _10458_ ;
wire _10459_ ;
wire _10460_ ;
wire _10461_ ;
wire _10462_ ;
wire _10463_ ;
wire _10464_ ;
wire _10465_ ;
wire _10466_ ;
wire _10467_ ;
wire _10468_ ;
wire _10469_ ;
wire _10470_ ;
wire _10471_ ;
wire _10472_ ;
wire _10473_ ;
wire _10474_ ;
wire _10475_ ;
wire _10476_ ;
wire _10477_ ;
wire _10478_ ;
wire _10479_ ;
wire _10480_ ;
wire _10481_ ;
wire _10482_ ;
wire _10483_ ;
wire _10484_ ;
wire _10485_ ;
wire _10486_ ;
wire _10487_ ;
wire _10488_ ;
wire _10489_ ;
wire _10490_ ;
wire _10491_ ;
wire _10492_ ;
wire _10493_ ;
wire _10494_ ;
wire _10495_ ;
wire _10496_ ;
wire _10497_ ;
wire _10498_ ;
wire _10499_ ;
wire _10500_ ;
wire _10501_ ;
wire _10502_ ;
wire _10503_ ;
wire _10504_ ;
wire _10505_ ;
wire _10506_ ;
wire _10507_ ;
wire _10508_ ;
wire _10509_ ;
wire _10510_ ;
wire _10511_ ;
wire _10512_ ;
wire _10513_ ;
wire _10514_ ;
wire _10515_ ;
wire _10516_ ;
wire _10517_ ;
wire _10518_ ;
wire _10519_ ;
wire _10520_ ;
wire _10521_ ;
wire _10522_ ;
wire _10523_ ;
wire _10524_ ;
wire _10525_ ;
wire _10526_ ;
wire _10527_ ;
wire _10528_ ;
wire _10529_ ;
wire _10530_ ;
wire _10531_ ;
wire _10532_ ;
wire _10533_ ;
wire _10534_ ;
wire _10535_ ;
wire _10536_ ;
wire _10537_ ;
wire _10538_ ;
wire _10539_ ;
wire _10540_ ;
wire _10541_ ;
wire _10542_ ;
wire _10543_ ;
wire _10544_ ;
wire _10545_ ;
wire _10546_ ;
wire _10547_ ;
wire _10548_ ;
wire _10549_ ;
wire _10550_ ;
wire _10551_ ;
wire _10552_ ;
wire _10553_ ;
wire _10554_ ;
wire _10555_ ;
wire _10556_ ;
wire _10557_ ;
wire _10558_ ;
wire _10559_ ;
wire _10560_ ;
wire _10561_ ;
wire _10562_ ;
wire _10563_ ;
wire _10564_ ;
wire _10565_ ;
wire _10566_ ;
wire _10567_ ;
wire _10568_ ;
wire _10569_ ;
wire _10570_ ;
wire _10571_ ;
wire _10572_ ;
wire _10573_ ;
wire _10574_ ;
wire _10575_ ;
wire _10576_ ;
wire _10577_ ;
wire _10578_ ;
wire _10579_ ;
wire _10580_ ;
wire _10581_ ;
wire _10582_ ;
wire _10583_ ;
wire _10584_ ;
wire _10585_ ;
wire _10586_ ;
wire _10587_ ;
wire _10588_ ;
wire _10589_ ;
wire _10590_ ;
wire _10591_ ;
wire _10592_ ;
wire _10593_ ;
wire _10594_ ;
wire _10595_ ;
wire _10596_ ;
wire _10597_ ;
wire _10598_ ;
wire _10599_ ;
wire _10600_ ;
wire _10601_ ;
wire _10602_ ;
wire _10603_ ;
wire _10604_ ;
wire _10605_ ;
wire _10606_ ;
wire _10607_ ;
wire _10608_ ;
wire _10609_ ;
wire _10610_ ;
wire _10611_ ;
wire _10612_ ;
wire _10613_ ;
wire _10614_ ;
wire _10615_ ;
wire _10616_ ;
wire _10617_ ;
wire _10618_ ;
wire _10619_ ;
wire _10620_ ;
wire _10621_ ;
wire _10622_ ;
wire _10623_ ;
wire _10624_ ;
wire _10625_ ;
wire _10626_ ;
wire _10627_ ;
wire _10628_ ;
wire _10629_ ;
wire _10630_ ;
wire _10631_ ;
wire _10632_ ;
wire _10633_ ;
wire _10634_ ;
wire _10635_ ;
wire _10636_ ;
wire _10637_ ;
wire _10638_ ;
wire _10639_ ;
wire _10640_ ;
wire _10641_ ;
wire _10642_ ;
wire _10643_ ;
wire _10644_ ;
wire _10645_ ;
wire _10646_ ;
wire _10647_ ;
wire _10648_ ;
wire _10649_ ;
wire _10650_ ;
wire _10651_ ;
wire _10652_ ;
wire _10653_ ;
wire _10654_ ;
wire _10655_ ;
wire _10656_ ;
wire _10657_ ;
wire _10658_ ;
wire _10659_ ;
wire _10660_ ;
wire _10661_ ;
wire _10662_ ;
wire _10663_ ;
wire _10664_ ;
wire _10665_ ;
wire _10666_ ;
wire _10667_ ;
wire _10668_ ;
wire _10669_ ;
wire _10670_ ;
wire _10671_ ;
wire _10672_ ;
wire _10673_ ;
wire _10674_ ;
wire _10675_ ;
wire _10676_ ;
wire _10677_ ;
wire _10678_ ;
wire _10679_ ;
wire _10680_ ;
wire _10681_ ;
wire _10682_ ;
wire _10683_ ;
wire _10684_ ;
wire _10685_ ;
wire _10686_ ;
wire _10687_ ;
wire _10688_ ;
wire _10689_ ;
wire _10690_ ;
wire _10691_ ;
wire _10692_ ;
wire _10693_ ;
wire _10694_ ;
wire _10695_ ;
wire _10696_ ;
wire _10697_ ;
wire _10698_ ;
wire _10699_ ;
wire _10700_ ;
wire _10701_ ;
wire _10702_ ;
wire _10703_ ;
wire _10704_ ;
wire _10705_ ;
wire _10706_ ;
wire _10707_ ;
wire _10708_ ;
wire _10709_ ;
wire _10710_ ;
wire _10711_ ;
wire _10712_ ;
wire _10713_ ;
wire _10714_ ;
wire _10715_ ;
wire _10716_ ;
wire _10717_ ;
wire _10718_ ;
wire _10719_ ;
wire _10720_ ;
wire _10721_ ;
wire _10722_ ;
wire _10723_ ;
wire _10724_ ;
wire _10725_ ;
wire _10726_ ;
wire _10727_ ;
wire _10728_ ;
wire _10729_ ;
wire _10730_ ;
wire _10731_ ;
wire _10732_ ;
wire _10733_ ;
wire _10734_ ;
wire _10735_ ;
wire _10736_ ;
wire _10737_ ;
wire _10738_ ;
wire _10739_ ;
wire _10740_ ;
wire _10741_ ;
wire _10742_ ;
wire _10743_ ;
wire _10744_ ;
wire _10745_ ;
wire _10746_ ;
wire _10747_ ;
wire _10748_ ;
wire _10749_ ;
wire _10750_ ;
wire _10751_ ;
wire _10752_ ;
wire _10753_ ;
wire _10754_ ;
wire _10755_ ;
wire _10756_ ;
wire _10757_ ;
wire _10758_ ;
wire _10759_ ;
wire _10760_ ;
wire _10761_ ;
wire _10762_ ;
wire _10763_ ;
wire _10764_ ;
wire _10765_ ;
wire _10766_ ;
wire _10767_ ;
wire _10768_ ;
wire _10769_ ;
wire _10770_ ;
wire _10771_ ;
wire _10772_ ;
wire _10773_ ;
wire _10774_ ;
wire _10775_ ;
wire _10776_ ;
wire _10777_ ;
wire _10778_ ;
wire _10779_ ;
wire _10780_ ;
wire _10781_ ;
wire _10782_ ;
wire _10783_ ;
wire _10784_ ;
wire _10785_ ;
wire _10786_ ;
wire _10787_ ;
wire _10788_ ;
wire _10789_ ;
wire _10790_ ;
wire _10791_ ;
wire _10792_ ;
wire _10793_ ;
wire _10794_ ;
wire _10795_ ;
wire _10796_ ;
wire _10797_ ;
wire _10798_ ;
wire _10799_ ;
wire _10800_ ;
wire _10801_ ;
wire _10802_ ;
wire _10803_ ;
wire _10804_ ;
wire _10805_ ;
wire _10806_ ;
wire _10807_ ;
wire _10808_ ;
wire _10809_ ;
wire _10810_ ;
wire _10811_ ;
wire _10812_ ;
wire _10813_ ;
wire _10814_ ;
wire _10815_ ;
wire _10816_ ;
wire _10817_ ;
wire _10818_ ;
wire _10819_ ;
wire _10820_ ;
wire _10821_ ;
wire _10822_ ;
wire _10823_ ;
wire _10824_ ;
wire _10825_ ;
wire _10826_ ;
wire _10827_ ;
wire _10828_ ;
wire _10829_ ;
wire _10830_ ;
wire _10831_ ;
wire _10832_ ;
wire _10833_ ;
wire _10834_ ;
wire _10835_ ;
wire _10836_ ;
wire _10837_ ;
wire _10838_ ;
wire _10839_ ;
wire _10840_ ;
wire _10841_ ;
wire _10842_ ;
wire _10843_ ;
wire _10844_ ;
wire _10845_ ;
wire _10846_ ;
wire _10847_ ;
wire _10848_ ;
wire _10849_ ;
wire _10850_ ;
wire _10851_ ;
wire _10852_ ;
wire _10853_ ;
wire _10854_ ;
wire _10855_ ;
wire _10856_ ;
wire _10857_ ;
wire _10858_ ;
wire _10859_ ;
wire _10860_ ;
wire _10861_ ;
wire _10862_ ;
wire _10863_ ;
wire _10864_ ;
wire _10865_ ;
wire _10866_ ;
wire _10867_ ;
wire _10868_ ;
wire _10869_ ;
wire _10870_ ;
wire _10871_ ;
wire _10872_ ;
wire _10873_ ;
wire _10874_ ;
wire _10875_ ;
wire _10876_ ;
wire _10877_ ;
wire _10878_ ;
wire _10879_ ;
wire _10880_ ;
wire _10881_ ;
wire _10882_ ;
wire _10883_ ;
wire _10884_ ;
wire _10885_ ;
wire _10886_ ;
wire _10887_ ;
wire _10888_ ;
wire _10889_ ;
wire _10890_ ;
wire _10891_ ;
wire _10892_ ;
wire _10893_ ;
wire _10894_ ;
wire _10895_ ;
wire _10896_ ;
wire _10897_ ;
wire _10898_ ;
wire _10899_ ;
wire _10900_ ;
wire _10901_ ;
wire _10902_ ;
wire _10903_ ;
wire _10904_ ;
wire _10905_ ;
wire _10906_ ;
wire _10907_ ;
wire _10908_ ;
wire _10909_ ;
wire _10910_ ;
wire _10911_ ;
wire _10912_ ;
wire _10913_ ;
wire _10914_ ;
wire _10915_ ;
wire _10916_ ;
wire _10917_ ;
wire _10918_ ;
wire _10919_ ;
wire _10920_ ;
wire _10921_ ;
wire _10922_ ;
wire _10923_ ;
wire _10924_ ;
wire _10925_ ;
wire _10926_ ;
wire _10927_ ;
wire _10928_ ;
wire _10929_ ;
wire _10930_ ;
wire _10931_ ;
wire _10932_ ;
wire _10933_ ;
wire _10934_ ;
wire _10935_ ;
wire _10936_ ;
wire _10937_ ;
wire _10938_ ;
wire _10939_ ;
wire _10940_ ;
wire _10941_ ;
wire _10942_ ;
wire _10943_ ;
wire _10944_ ;
wire _10945_ ;
wire _10946_ ;
wire _10947_ ;
wire _10948_ ;
wire _10949_ ;
wire _10950_ ;
wire _10951_ ;
wire _10952_ ;
wire _10953_ ;
wire _10954_ ;
wire _10955_ ;
wire _10956_ ;
wire _10957_ ;
wire _10958_ ;
wire _10959_ ;
wire _10960_ ;
wire _10961_ ;
wire _10962_ ;
wire _10963_ ;
wire _10964_ ;
wire _10965_ ;
wire _10966_ ;
wire _10967_ ;
wire _10968_ ;
wire _10969_ ;
wire _10970_ ;
wire _10971_ ;
wire _10972_ ;
wire _10973_ ;
wire _10974_ ;
wire _10975_ ;
wire _10976_ ;
wire _10977_ ;
wire _10978_ ;
wire _10979_ ;
wire _10980_ ;
wire _10981_ ;
wire _10982_ ;
wire _10983_ ;
wire _10984_ ;
wire _10985_ ;
wire _10986_ ;
wire _10987_ ;
wire _10988_ ;
wire _10989_ ;
wire _10990_ ;
wire _10991_ ;
wire _10992_ ;
wire _10993_ ;
wire _10994_ ;
wire _10995_ ;
wire _10996_ ;
wire _10997_ ;
wire _10998_ ;
wire _10999_ ;
wire _11000_ ;
wire _11001_ ;
wire _11002_ ;
wire _11003_ ;
wire _11004_ ;
wire _11005_ ;
wire _11006_ ;
wire _11007_ ;
wire _11008_ ;
wire _11009_ ;
wire _11010_ ;
wire _11011_ ;
wire _11012_ ;
wire _11013_ ;
wire _11014_ ;
wire _11015_ ;
wire _11016_ ;
wire _11017_ ;
wire _11018_ ;
wire _11019_ ;
wire _11020_ ;
wire _11021_ ;
wire _11022_ ;
wire _11023_ ;
wire _11024_ ;
wire _11025_ ;
wire _11026_ ;
wire _11027_ ;
wire _11028_ ;
wire _11029_ ;
wire _11030_ ;
wire _11031_ ;
wire _11032_ ;
wire _11033_ ;
wire _11034_ ;
wire _11035_ ;
wire _11036_ ;
wire _11037_ ;
wire _11038_ ;
wire _11039_ ;
wire _11040_ ;
wire _11041_ ;
wire _11042_ ;
wire _11043_ ;
wire _11044_ ;
wire _11045_ ;
wire _11046_ ;
wire _11047_ ;
wire _11048_ ;
wire _11049_ ;
wire _11050_ ;
wire _11051_ ;
wire _11052_ ;
wire _11053_ ;
wire _11054_ ;
wire _11055_ ;
wire _11056_ ;
wire _11057_ ;
wire _11058_ ;
wire _11059_ ;
wire _11060_ ;
wire _11061_ ;
wire _11062_ ;
wire _11063_ ;
wire _11064_ ;
wire _11065_ ;
wire _11066_ ;
wire _11067_ ;
wire _11068_ ;
wire _11069_ ;
wire _11070_ ;
wire _11071_ ;
wire _11072_ ;
wire _11073_ ;
wire _11074_ ;
wire _11075_ ;
wire _11076_ ;
wire _11077_ ;
wire _11078_ ;
wire _11079_ ;
wire _11080_ ;
wire _11081_ ;
wire _11082_ ;
wire _11083_ ;
wire _11084_ ;
wire _11085_ ;
wire _11086_ ;
wire _11087_ ;
wire _11088_ ;
wire _11089_ ;
wire _11090_ ;
wire _11091_ ;
wire _11092_ ;
wire _11093_ ;
wire _11094_ ;
wire _11095_ ;
wire _11096_ ;
wire _11097_ ;
wire _11098_ ;
wire _11099_ ;
wire _11100_ ;
wire _11101_ ;
wire _11102_ ;
wire _11103_ ;
wire _11104_ ;
wire _11105_ ;
wire _11106_ ;
wire _11107_ ;
wire _11108_ ;
wire _11109_ ;
wire _11110_ ;
wire _11111_ ;
wire _11112_ ;
wire _11113_ ;
wire _11114_ ;
wire _11115_ ;
wire _11116_ ;
wire _11117_ ;
wire _11118_ ;
wire _11119_ ;
wire _11120_ ;
wire _11121_ ;
wire _11122_ ;
wire _11123_ ;
wire _11124_ ;
wire _11125_ ;
wire _11126_ ;
wire _11127_ ;
wire _11128_ ;
wire _11129_ ;
wire _11130_ ;
wire _11131_ ;
wire _11132_ ;
wire _11133_ ;
wire _11134_ ;
wire _11135_ ;
wire _11136_ ;
wire _11137_ ;
wire _11138_ ;
wire _11139_ ;
wire _11140_ ;
wire _11141_ ;
wire _11142_ ;
wire _11143_ ;
wire _11144_ ;
wire _11145_ ;
wire _11146_ ;
wire _11147_ ;
wire _11148_ ;
wire _11149_ ;
wire _11150_ ;
wire _11151_ ;
wire _11152_ ;
wire _11153_ ;
wire _11154_ ;
wire _11155_ ;
wire _11156_ ;
wire _11157_ ;
wire _11158_ ;
wire _11159_ ;
wire _11160_ ;
wire _11161_ ;
wire _11162_ ;
wire _11163_ ;
wire _11164_ ;
wire _11165_ ;
wire _11166_ ;
wire _11167_ ;
wire _11168_ ;
wire _11169_ ;
wire _11170_ ;
wire _11171_ ;
wire _11172_ ;
wire _11173_ ;
wire _11174_ ;
wire _11175_ ;
wire _11176_ ;
wire _11177_ ;
wire _11178_ ;
wire _11179_ ;
wire _11180_ ;
wire _11181_ ;
wire _11182_ ;
wire _11183_ ;
wire _11184_ ;
wire _11185_ ;
wire _11186_ ;
wire _11187_ ;
wire _11188_ ;
wire _11189_ ;
wire _11190_ ;
wire _11191_ ;
wire _11192_ ;
wire _11193_ ;
wire _11194_ ;
wire _11195_ ;
wire _11196_ ;
wire _11197_ ;
wire _11198_ ;
wire _11199_ ;
wire _11200_ ;
wire _11201_ ;
wire _11202_ ;
wire _11203_ ;
wire _11204_ ;
wire _11205_ ;
wire _11206_ ;
wire _11207_ ;
wire _11208_ ;
wire _11209_ ;
wire _11210_ ;
wire _11211_ ;
wire _11212_ ;
wire _11213_ ;
wire _11214_ ;
wire _11215_ ;
wire _11216_ ;
wire _11217_ ;
wire _11218_ ;
wire _11219_ ;
wire _11220_ ;
wire _11221_ ;
wire _11222_ ;
wire _11223_ ;
wire _11224_ ;
wire _11225_ ;
wire _11226_ ;
wire _11227_ ;
wire _11228_ ;
wire _11229_ ;
wire _11230_ ;
wire _11231_ ;
wire _11232_ ;
wire _11233_ ;
wire _11234_ ;
wire _11235_ ;
wire _11236_ ;
wire _11237_ ;
wire _11238_ ;
wire _11239_ ;
wire _11240_ ;
wire _11241_ ;
wire _11242_ ;
wire _11243_ ;
wire _11244_ ;
wire _11245_ ;
wire _11246_ ;
wire _11247_ ;
wire _11248_ ;
wire _11249_ ;
wire _11250_ ;
wire _11251_ ;
wire _11252_ ;
wire _11253_ ;
wire _11254_ ;
wire _11255_ ;
wire _11256_ ;
wire _11257_ ;
wire _11258_ ;
wire _11259_ ;
wire _11260_ ;
wire _11261_ ;
wire _11262_ ;
wire _11263_ ;
wire _11264_ ;
wire _11265_ ;
wire _11266_ ;
wire _11267_ ;
wire _11268_ ;
wire _11269_ ;
wire _11270_ ;
wire _11271_ ;
wire _11272_ ;
wire _11273_ ;
wire _11274_ ;
wire _11275_ ;
wire _11276_ ;
wire _11277_ ;
wire _11278_ ;
wire _11279_ ;
wire _11280_ ;
wire _11281_ ;
wire _11282_ ;
wire _11283_ ;
wire _11284_ ;
wire _11285_ ;
wire _11286_ ;
wire _11287_ ;
wire _11288_ ;
wire _11289_ ;
wire _11290_ ;
wire _11291_ ;
wire _11292_ ;
wire _11293_ ;
wire _11294_ ;
wire _11295_ ;
wire _11296_ ;
wire _11297_ ;
wire _11298_ ;
wire _11299_ ;
wire _11300_ ;
wire _11301_ ;
wire _11302_ ;
wire _11303_ ;
wire _11304_ ;
wire _11305_ ;
wire _11306_ ;
wire _11307_ ;
wire _11308_ ;
wire _11309_ ;
wire _11310_ ;
wire _11311_ ;
wire _11312_ ;
wire _11313_ ;
wire _11314_ ;
wire _11315_ ;
wire _11316_ ;
wire _11317_ ;
wire _11318_ ;
wire _11319_ ;
wire _11320_ ;
wire _11321_ ;
wire _11322_ ;
wire _11323_ ;
wire _11324_ ;
wire _11325_ ;
wire _11326_ ;
wire _11327_ ;
wire _11328_ ;
wire _11329_ ;
wire _11330_ ;
wire _11331_ ;
wire _11332_ ;
wire _11333_ ;
wire _11334_ ;
wire _11335_ ;
wire _11336_ ;
wire _11337_ ;
wire _11338_ ;
wire _11339_ ;
wire _11340_ ;
wire _11341_ ;
wire _11342_ ;
wire _11343_ ;
wire _11344_ ;
wire _11345_ ;
wire _11346_ ;
wire _11347_ ;
wire _11348_ ;
wire _11349_ ;
wire _11350_ ;
wire _11351_ ;
wire _11352_ ;
wire _11353_ ;
wire _11354_ ;
wire _11355_ ;
wire _11356_ ;
wire _11357_ ;
wire _11358_ ;
wire _11359_ ;
wire _11360_ ;
wire _11361_ ;
wire _11362_ ;
wire _11363_ ;
wire _11364_ ;
wire _11365_ ;
wire _11366_ ;
wire _11367_ ;
wire _11368_ ;
wire _11369_ ;
wire _11370_ ;
wire _11371_ ;
wire _11372_ ;
wire _11373_ ;
wire _11374_ ;
wire _11375_ ;
wire _11376_ ;
wire _11377_ ;
wire _11378_ ;
wire _11379_ ;
wire _11380_ ;
wire _11381_ ;
wire _11382_ ;
wire _11383_ ;
wire _11384_ ;
wire _11385_ ;
wire _11386_ ;
wire _11387_ ;
wire _11388_ ;
wire _11389_ ;
wire _11390_ ;
wire _11391_ ;
wire _11392_ ;
wire _11393_ ;
wire _11394_ ;
wire _11395_ ;
wire _11396_ ;
wire _11397_ ;
wire _11398_ ;
wire _11399_ ;
wire _11400_ ;
wire _11401_ ;
wire _11402_ ;
wire _11403_ ;
wire _11404_ ;
wire _11405_ ;
wire _11406_ ;
wire _11407_ ;
wire _11408_ ;
wire _11409_ ;
wire _11410_ ;
wire _11411_ ;
wire _11412_ ;
wire _11413_ ;
wire _11414_ ;
wire _11415_ ;
wire _11416_ ;
wire _11417_ ;
wire _11418_ ;
wire _11419_ ;
wire _11420_ ;
wire _11421_ ;
wire _11422_ ;
wire _11423_ ;
wire _11424_ ;
wire _11425_ ;
wire _11426_ ;
wire _11427_ ;
wire _11428_ ;
wire _11429_ ;
wire _11430_ ;
wire _11431_ ;
wire _11432_ ;
wire _11433_ ;
wire _11434_ ;
wire _11435_ ;
wire _11436_ ;
wire _11437_ ;
wire _11438_ ;
wire _11439_ ;
wire _11440_ ;
wire _11441_ ;
wire _11442_ ;
wire _11443_ ;
wire _11444_ ;
wire _11445_ ;
wire _11446_ ;
wire _11447_ ;
wire _11448_ ;
wire _11449_ ;
wire _11450_ ;
wire _11451_ ;
wire _11452_ ;
wire _11453_ ;
wire _11454_ ;
wire _11455_ ;
wire _11456_ ;
wire _11457_ ;
wire _11458_ ;
wire _11459_ ;
wire _11460_ ;
wire _11461_ ;
wire _11462_ ;
wire _11463_ ;
wire _11464_ ;
wire _11465_ ;
wire _11466_ ;
wire _11467_ ;
wire _11468_ ;
wire _11469_ ;
wire _11470_ ;
wire _11471_ ;
wire _11472_ ;
wire _11473_ ;
wire _11474_ ;
wire _11475_ ;
wire _11476_ ;
wire _11477_ ;
wire _11478_ ;
wire _11479_ ;
wire _11480_ ;
wire _11481_ ;
wire _11482_ ;
wire _11483_ ;
wire _11484_ ;
wire _11485_ ;
wire _11486_ ;
wire _11487_ ;
wire _11488_ ;
wire _11489_ ;
wire _11490_ ;
wire _11491_ ;
wire _11492_ ;
wire _11493_ ;
wire _11494_ ;
wire _11495_ ;
wire _11496_ ;
wire _11497_ ;
wire _11498_ ;
wire _11499_ ;
wire _11500_ ;
wire _11501_ ;
wire _11502_ ;
wire _11503_ ;
wire _11504_ ;
wire _11505_ ;
wire _11506_ ;
wire _11507_ ;
wire _11508_ ;
wire _11509_ ;
wire _11510_ ;
wire _11511_ ;
wire _11512_ ;
wire _11513_ ;
wire _11514_ ;
wire _11515_ ;
wire _11516_ ;
wire _11517_ ;
wire _11518_ ;
wire _11519_ ;
wire _11520_ ;
wire _11521_ ;
wire _11522_ ;
wire _11523_ ;
wire _11524_ ;
wire _11525_ ;
wire _11526_ ;
wire _11527_ ;
wire _11528_ ;
wire _11529_ ;
wire _11530_ ;
wire _11531_ ;
wire _11532_ ;
wire _11533_ ;
wire _11534_ ;
wire _11535_ ;
wire _11536_ ;
wire _11537_ ;
wire _11538_ ;
wire _11539_ ;
wire _11540_ ;
wire _11541_ ;
wire _11542_ ;
wire _11543_ ;
wire _11544_ ;
wire _11545_ ;
wire _11546_ ;
wire _11547_ ;
wire _11548_ ;
wire _11549_ ;
wire _11550_ ;
wire _11551_ ;
wire _11552_ ;
wire _11553_ ;
wire _11554_ ;
wire _11555_ ;
wire _11556_ ;
wire _11557_ ;
wire _11558_ ;
wire _11559_ ;
wire _11560_ ;
wire _11561_ ;
wire _11562_ ;
wire _11563_ ;
wire _11564_ ;
wire _11565_ ;
wire _11566_ ;
wire _11567_ ;
wire _11568_ ;
wire _11569_ ;
wire _11570_ ;
wire _11571_ ;
wire _11572_ ;
wire _11573_ ;
wire _11574_ ;
wire _11575_ ;
wire _11576_ ;
wire _11577_ ;
wire _11578_ ;
wire _11579_ ;
wire _11580_ ;
wire _11581_ ;
wire _11582_ ;
wire _11583_ ;
wire _11584_ ;
wire _11585_ ;
wire _11586_ ;
wire _11587_ ;
wire _11588_ ;
wire _11589_ ;
wire _11590_ ;
wire _11591_ ;
wire _11592_ ;
wire _11593_ ;
wire _11594_ ;
wire _11595_ ;
wire _11596_ ;
wire _11597_ ;
wire _11598_ ;
wire _11599_ ;
wire _11600_ ;
wire _11601_ ;
wire _11602_ ;
wire _11603_ ;
wire _11604_ ;
wire _11605_ ;
wire _11606_ ;
wire _11607_ ;
wire _11608_ ;
wire _11609_ ;
wire _11610_ ;
wire _11611_ ;
wire _11612_ ;
wire _11613_ ;
wire _11614_ ;
wire _11615_ ;
wire _11616_ ;
wire _11617_ ;
wire _11618_ ;
wire _11619_ ;
wire _11620_ ;
wire _11621_ ;
wire _11622_ ;
wire _11623_ ;
wire _11624_ ;
wire _11625_ ;
wire _11626_ ;
wire _11627_ ;
wire _11628_ ;
wire _11629_ ;
wire _11630_ ;
wire _11631_ ;
wire _11632_ ;
wire _11633_ ;
wire _11634_ ;
wire _11635_ ;
wire _11636_ ;
wire _11637_ ;
wire _11638_ ;
wire _11639_ ;
wire _11640_ ;
wire _11641_ ;
wire _11642_ ;
wire _11643_ ;
wire _11644_ ;
wire _11645_ ;
wire _11646_ ;
wire _11647_ ;
wire _11648_ ;
wire _11649_ ;
wire _11650_ ;
wire _11651_ ;
wire _11652_ ;
wire _11653_ ;
wire _11654_ ;
wire _11655_ ;
wire _11656_ ;
wire _11657_ ;
wire _11658_ ;
wire _11659_ ;
wire _11660_ ;
wire _11661_ ;
wire _11662_ ;
wire _11663_ ;
wire _11664_ ;
wire _11665_ ;
wire _11666_ ;
wire _11667_ ;
wire _11668_ ;
wire _11669_ ;
wire _11670_ ;
wire _11671_ ;
wire _11672_ ;
wire _11673_ ;
wire _11674_ ;
wire _11675_ ;
wire _11676_ ;
wire _11677_ ;
wire _11678_ ;
wire _11679_ ;
wire _11680_ ;
wire _11681_ ;
wire _11682_ ;
wire _11683_ ;
wire _11684_ ;
wire _11685_ ;
wire _11686_ ;
wire _11687_ ;
wire _11688_ ;
wire _11689_ ;
wire _11690_ ;
wire _11691_ ;
wire _11692_ ;
wire _11693_ ;
wire _11694_ ;
wire _11695_ ;
wire _11696_ ;
wire _11697_ ;
wire _11698_ ;
wire _11699_ ;
wire _11700_ ;
wire _11701_ ;
wire _11702_ ;
wire _11703_ ;
wire _11704_ ;
wire _11705_ ;
wire _11706_ ;
wire _11707_ ;
wire _11708_ ;
wire _11709_ ;
wire _11710_ ;
wire _11711_ ;
wire _11712_ ;
wire _11713_ ;
wire _11714_ ;
wire _11715_ ;
wire _11716_ ;
wire _11717_ ;
wire _11718_ ;
wire _11719_ ;
wire _11720_ ;
wire _11721_ ;
wire _11722_ ;
wire _11723_ ;
wire _11724_ ;
wire _11725_ ;
wire _11726_ ;
wire _11727_ ;
wire _11728_ ;
wire _11729_ ;
wire _11730_ ;
wire _11731_ ;
wire _11732_ ;
wire _11733_ ;
wire _11734_ ;
wire _11735_ ;
wire _11736_ ;
wire _11737_ ;
wire _11738_ ;
wire _11739_ ;
wire _11740_ ;
wire _11741_ ;
wire _11742_ ;
wire _11743_ ;
wire _11744_ ;
wire _11745_ ;
wire _11746_ ;
wire _11747_ ;
wire _11748_ ;
wire _11749_ ;
wire _11750_ ;
wire _11751_ ;
wire _11752_ ;
wire _11753_ ;
wire _11754_ ;
wire _11755_ ;
wire _11756_ ;
wire _11757_ ;
wire _11758_ ;
wire _11759_ ;
wire _11760_ ;
wire _11761_ ;
wire _11762_ ;
wire _11763_ ;
wire _11764_ ;
wire _11765_ ;
wire _11766_ ;
wire _11767_ ;
wire _11768_ ;
wire _11769_ ;
wire _11770_ ;
wire _11771_ ;
wire _11772_ ;
wire _11773_ ;
wire _11774_ ;
wire _11775_ ;
wire _11776_ ;
wire _11777_ ;
wire _11778_ ;
wire _11779_ ;
wire _11780_ ;
wire _11781_ ;
wire _11782_ ;
wire _11783_ ;
wire _11784_ ;
wire _11785_ ;
wire _11786_ ;
wire _11787_ ;
wire _11788_ ;
wire _11789_ ;
wire _11790_ ;
wire _11791_ ;
wire _11792_ ;
wire _11793_ ;
wire _11794_ ;
wire _11795_ ;
wire _11796_ ;
wire _11797_ ;
wire _11798_ ;
wire _11799_ ;
wire _11800_ ;
wire _11801_ ;
wire _11802_ ;
wire _11803_ ;
wire _11804_ ;
wire _11805_ ;
wire _11806_ ;
wire _11807_ ;
wire _11808_ ;
wire _11809_ ;
wire _11810_ ;
wire _11811_ ;
wire _11812_ ;
wire _11813_ ;
wire _11814_ ;
wire _11815_ ;
wire _11816_ ;
wire _11817_ ;
wire _11818_ ;
wire _11819_ ;
wire _11820_ ;
wire _11821_ ;
wire _11822_ ;
wire _11823_ ;
wire _11824_ ;
wire _11825_ ;
wire _11826_ ;
wire _11827_ ;
wire _11828_ ;
wire _11829_ ;
wire _11830_ ;
wire _11831_ ;
wire _11832_ ;
wire _11833_ ;
wire _11834_ ;
wire _11835_ ;
wire _11836_ ;
wire _11837_ ;
wire _11838_ ;
wire _11839_ ;
wire _11840_ ;
wire _11841_ ;
wire _11842_ ;
wire _11843_ ;
wire _11844_ ;
wire _11845_ ;
wire _11846_ ;
wire _11847_ ;
wire _11848_ ;
wire _11849_ ;
wire _11850_ ;
wire _11851_ ;
wire _11852_ ;
wire _11853_ ;
wire _11854_ ;
wire _11855_ ;
wire _11856_ ;
wire _11857_ ;
wire _11858_ ;
wire _11859_ ;
wire _11860_ ;
wire _11861_ ;
wire _11862_ ;
wire _11863_ ;
wire _11864_ ;
wire _11865_ ;
wire _11866_ ;
wire _11867_ ;
wire _11868_ ;
wire _11869_ ;
wire _11870_ ;
wire _11871_ ;
wire _11872_ ;
wire _11873_ ;
wire _11874_ ;
wire _11875_ ;
wire _11876_ ;
wire _11877_ ;
wire _11878_ ;
wire _11879_ ;
wire _11880_ ;
wire _11881_ ;
wire _11882_ ;
wire _11883_ ;
wire _11884_ ;
wire _11885_ ;
wire _11886_ ;
wire _11887_ ;
wire _11888_ ;
wire _11889_ ;
wire _11890_ ;
wire _11891_ ;
wire _11892_ ;
wire _11893_ ;
wire _11894_ ;
wire _11895_ ;
wire _11896_ ;
wire _11897_ ;
wire _11898_ ;
wire _11899_ ;
wire _11900_ ;
wire _11901_ ;
wire _11902_ ;
wire _11903_ ;
wire _11904_ ;
wire _11905_ ;
wire _11906_ ;
wire _11907_ ;
wire _11908_ ;
wire _11909_ ;
wire _11910_ ;
wire _11911_ ;
wire _11912_ ;
wire _11913_ ;
wire _11914_ ;
wire _11915_ ;
wire _11916_ ;
wire _11917_ ;
wire _11918_ ;
wire _11919_ ;
wire _11920_ ;
wire _11921_ ;
wire _11922_ ;
wire _11923_ ;
wire _11924_ ;
wire _11925_ ;
wire _11926_ ;
wire _11927_ ;
wire _11928_ ;
wire _11929_ ;
wire _11930_ ;
wire _11931_ ;
wire _11932_ ;
wire _11933_ ;
wire _11934_ ;
wire _11935_ ;
wire _11936_ ;
wire _11937_ ;
wire _11938_ ;
wire _11939_ ;
wire _11940_ ;
wire _11941_ ;
wire _11942_ ;
wire _11943_ ;
wire _11944_ ;
wire _11945_ ;
wire _11946_ ;
wire _11947_ ;
wire _11948_ ;
wire _11949_ ;
wire _11950_ ;
wire _11951_ ;
wire _11952_ ;
wire _11953_ ;
wire _11954_ ;
wire _11955_ ;
wire _11956_ ;
wire _11957_ ;
wire _11958_ ;
wire _11959_ ;
wire _11960_ ;
wire _11961_ ;
wire _11962_ ;
wire _11963_ ;
wire _11964_ ;
wire _11965_ ;
wire _11966_ ;
wire _11967_ ;
wire _11968_ ;
wire _11969_ ;
wire _11970_ ;
wire _11971_ ;
wire _11972_ ;
wire _11973_ ;
wire _11974_ ;
wire _11975_ ;
wire _11976_ ;
wire _11977_ ;
wire _11978_ ;
wire _11979_ ;
wire _11980_ ;
wire _11981_ ;
wire _11982_ ;
wire _11983_ ;
wire _11984_ ;
wire _11985_ ;
wire _11986_ ;
wire _11987_ ;
wire _11988_ ;
wire _11989_ ;
wire _11990_ ;
wire _11991_ ;
wire _11992_ ;
wire _11993_ ;
wire _11994_ ;
wire _11995_ ;
wire _11996_ ;
wire _11997_ ;
wire _11998_ ;
wire _11999_ ;
wire _12000_ ;
wire _12001_ ;
wire _12002_ ;
wire _12003_ ;
wire _12004_ ;
wire _12005_ ;
wire _12006_ ;
wire _12007_ ;
wire _12008_ ;
wire _12009_ ;
wire _12010_ ;
wire _12011_ ;
wire _12012_ ;
wire _12013_ ;
wire _12014_ ;
wire _12015_ ;
wire _12016_ ;
wire _12017_ ;
wire _12018_ ;
wire _12019_ ;
wire _12020_ ;
wire _12021_ ;
wire alu_result_out_$_XNOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B_$_ORNOT__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B ;
wire alu_result_out_$_XNOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B_$_OR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire alu_result_out_$_XNOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__B_Y ;
wire alu_result_out_$_XNOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B_$_OR__Y_B_$_NOR__Y_A_$_XOR__Y_B_$_OR__Y_A_$_OR__Y_B ;
wire clk ;
wire dnpc_$_MUX__Y_11_A_$_NOT__Y_A_$_XOR__Y_B ;
wire dnpc_$_MUX__Y_13_A_$_NOT__Y_A_$_XOR__Y_B ;
wire dnpc_$_MUX__Y_15_A_$_NOT__Y_A_$_XOR__Y_B ;
wire dnpc_$_MUX__Y_17_A_$_NOT__Y_A_$_XOR__Y_B ;
wire dnpc_$_MUX__Y_1_A_$_NOT__Y_A_$_XOR__Y_B ;
wire dnpc_$_MUX__Y_21_A_$_NOT__Y_A_$_XOR__Y_B ;
wire dnpc_$_MUX__Y_22_A ;
wire dnpc_$_MUX__Y_3_A_$_NOT__Y_A_$_XOR__Y_B ;
wire dnpc_$_MUX__Y_5_A_$_NOT__Y_A_$_XOR__Y_B ;
wire dnpc_$_MUX__Y_9_A_$_NOT__Y_A_$_XOR__Y_B ;
wire dnpc_$_NOT__Y_1_A_$_MUX__Y_A_$_XOR__Y_B ;
wire dnpc_$_NOT__Y_3_A_$_MUX__Y_A_$_XOR__Y_B ;
wire dnpc_$_NOT__Y_5_A_$_MUX__Y_A_$_XOR__Y_B ;
wire dnpc_$_NOT__Y_A_$_ANDNOT__B_A ;
wire jump_en ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire reset ;
wire \u_gpr.gpr_wdata_$_ANDNOT__Y_30_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \u_gpr.regfile[0][0] ;
wire \u_gpr.regfile[0][10] ;
wire \u_gpr.regfile[0][11] ;
wire \u_gpr.regfile[0][12] ;
wire \u_gpr.regfile[0][13] ;
wire \u_gpr.regfile[0][14] ;
wire \u_gpr.regfile[0][15] ;
wire \u_gpr.regfile[0][16] ;
wire \u_gpr.regfile[0][17] ;
wire \u_gpr.regfile[0][18] ;
wire \u_gpr.regfile[0][19] ;
wire \u_gpr.regfile[0][1] ;
wire \u_gpr.regfile[0][20] ;
wire \u_gpr.regfile[0][21] ;
wire \u_gpr.regfile[0][22] ;
wire \u_gpr.regfile[0][23] ;
wire \u_gpr.regfile[0][24] ;
wire \u_gpr.regfile[0][25] ;
wire \u_gpr.regfile[0][26] ;
wire \u_gpr.regfile[0][27] ;
wire \u_gpr.regfile[0][28] ;
wire \u_gpr.regfile[0][29] ;
wire \u_gpr.regfile[0][2] ;
wire \u_gpr.regfile[0][30] ;
wire \u_gpr.regfile[0][31] ;
wire \u_gpr.regfile[0][3] ;
wire \u_gpr.regfile[0][4] ;
wire \u_gpr.regfile[0][5] ;
wire \u_gpr.regfile[0][6] ;
wire \u_gpr.regfile[0][7] ;
wire \u_gpr.regfile[0][8] ;
wire \u_gpr.regfile[0][9] ;
wire \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_E ;
wire \u_gpr.regfile[1][0] ;
wire \u_gpr.regfile[1][10] ;
wire \u_gpr.regfile[1][11] ;
wire \u_gpr.regfile[1][12] ;
wire \u_gpr.regfile[1][13] ;
wire \u_gpr.regfile[1][14] ;
wire \u_gpr.regfile[1][15] ;
wire \u_gpr.regfile[1][16] ;
wire \u_gpr.regfile[1][17] ;
wire \u_gpr.regfile[1][18] ;
wire \u_gpr.regfile[1][19] ;
wire \u_gpr.regfile[1][1] ;
wire \u_gpr.regfile[1][20] ;
wire \u_gpr.regfile[1][21] ;
wire \u_gpr.regfile[1][22] ;
wire \u_gpr.regfile[1][23] ;
wire \u_gpr.regfile[1][24] ;
wire \u_gpr.regfile[1][25] ;
wire \u_gpr.regfile[1][26] ;
wire \u_gpr.regfile[1][27] ;
wire \u_gpr.regfile[1][28] ;
wire \u_gpr.regfile[1][29] ;
wire \u_gpr.regfile[1][2] ;
wire \u_gpr.regfile[1][30] ;
wire \u_gpr.regfile[1][31] ;
wire \u_gpr.regfile[1][3] ;
wire \u_gpr.regfile[1][4] ;
wire \u_gpr.regfile[1][5] ;
wire \u_gpr.regfile[1][6] ;
wire \u_gpr.regfile[1][7] ;
wire \u_gpr.regfile[1][8] ;
wire \u_gpr.regfile[1][9] ;
wire \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_E ;
wire \u_gpr.regfile[2][0] ;
wire \u_gpr.regfile[2][10] ;
wire \u_gpr.regfile[2][11] ;
wire \u_gpr.regfile[2][12] ;
wire \u_gpr.regfile[2][13] ;
wire \u_gpr.regfile[2][14] ;
wire \u_gpr.regfile[2][15] ;
wire \u_gpr.regfile[2][16] ;
wire \u_gpr.regfile[2][17] ;
wire \u_gpr.regfile[2][18] ;
wire \u_gpr.regfile[2][19] ;
wire \u_gpr.regfile[2][1] ;
wire \u_gpr.regfile[2][20] ;
wire \u_gpr.regfile[2][21] ;
wire \u_gpr.regfile[2][22] ;
wire \u_gpr.regfile[2][23] ;
wire \u_gpr.regfile[2][24] ;
wire \u_gpr.regfile[2][25] ;
wire \u_gpr.regfile[2][26] ;
wire \u_gpr.regfile[2][27] ;
wire \u_gpr.regfile[2][28] ;
wire \u_gpr.regfile[2][29] ;
wire \u_gpr.regfile[2][2] ;
wire \u_gpr.regfile[2][30] ;
wire \u_gpr.regfile[2][31] ;
wire \u_gpr.regfile[2][3] ;
wire \u_gpr.regfile[2][4] ;
wire \u_gpr.regfile[2][5] ;
wire \u_gpr.regfile[2][6] ;
wire \u_gpr.regfile[2][7] ;
wire \u_gpr.regfile[2][8] ;
wire \u_gpr.regfile[2][9] ;
wire \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_E ;
wire \u_gpr.regfile[3][0] ;
wire \u_gpr.regfile[3][10] ;
wire \u_gpr.regfile[3][11] ;
wire \u_gpr.regfile[3][12] ;
wire \u_gpr.regfile[3][13] ;
wire \u_gpr.regfile[3][14] ;
wire \u_gpr.regfile[3][15] ;
wire \u_gpr.regfile[3][16] ;
wire \u_gpr.regfile[3][17] ;
wire \u_gpr.regfile[3][18] ;
wire \u_gpr.regfile[3][19] ;
wire \u_gpr.regfile[3][1] ;
wire \u_gpr.regfile[3][20] ;
wire \u_gpr.regfile[3][21] ;
wire \u_gpr.regfile[3][22] ;
wire \u_gpr.regfile[3][23] ;
wire \u_gpr.regfile[3][24] ;
wire \u_gpr.regfile[3][25] ;
wire \u_gpr.regfile[3][26] ;
wire \u_gpr.regfile[3][27] ;
wire \u_gpr.regfile[3][28] ;
wire \u_gpr.regfile[3][29] ;
wire \u_gpr.regfile[3][2] ;
wire \u_gpr.regfile[3][30] ;
wire \u_gpr.regfile[3][31] ;
wire \u_gpr.regfile[3][3] ;
wire \u_gpr.regfile[3][4] ;
wire \u_gpr.regfile[3][5] ;
wire \u_gpr.regfile[3][6] ;
wire \u_gpr.regfile[3][7] ;
wire \u_gpr.regfile[3][8] ;
wire \u_gpr.regfile[3][9] ;
wire \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_E ;
wire \u_ifu.jump_en_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_NOR__Y_A_$_OR__Y_B ;
wire \u_ifu.reset_sync ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_6 ;
wire fanout_net_7 ;
wire fanout_net_8 ;
wire fanout_net_9 ;
wire fanout_net_10 ;
wire fanout_net_11 ;
wire fanout_net_12 ;
wire fanout_net_13 ;
wire fanout_net_14 ;
wire fanout_net_15 ;
wire fanout_net_16 ;
wire fanout_net_17 ;
wire fanout_net_18 ;
wire fanout_net_19 ;
wire fanout_net_20 ;
wire fanout_net_21 ;
wire fanout_net_22 ;
wire fanout_net_23 ;
wire fanout_net_24 ;
wire fanout_net_25 ;
wire fanout_net_26 ;
wire fanout_net_27 ;
wire fanout_net_28 ;
wire fanout_net_29 ;
wire fanout_net_30 ;
wire fanout_net_31 ;
wire fanout_net_32 ;
wire fanout_net_33 ;
wire fanout_net_34 ;
wire fanout_net_35 ;
wire fanout_net_36 ;
wire fanout_net_37 ;
wire fanout_net_38 ;
wire fanout_net_39 ;
wire fanout_net_40 ;
wire fanout_net_41 ;
wire fanout_net_42 ;
wire fanout_net_43 ;
wire fanout_net_44 ;
wire fanout_net_45 ;
wire fanout_net_46 ;
wire fanout_net_47 ;
wire fanout_net_48 ;
wire fanout_net_49 ;
wire fanout_net_50 ;
wire fanout_net_51 ;
wire fanout_net_52 ;
wire fanout_net_53 ;
wire fanout_net_54 ;
wire fanout_net_55 ;
wire fanout_net_56 ;
wire fanout_net_57 ;
wire fanout_net_58 ;
wire fanout_net_59 ;
wire fanout_net_60 ;
wire fanout_net_61 ;
wire fanout_net_62 ;
wire fanout_net_63 ;
wire fanout_net_64 ;
wire fanout_net_65 ;
wire fanout_net_66 ;
wire fanout_net_67 ;
wire fanout_net_68 ;
wire fanout_net_69 ;
wire fanout_net_70 ;
wire fanout_net_71 ;
wire fanout_net_72 ;
wire fanout_net_73 ;
wire fanout_net_74 ;
wire fanout_net_75 ;
wire fanout_net_76 ;
wire \alu_result_out[0] ;
wire \alu_result_out[1] ;
wire \alu_result_out[2] ;
wire \alu_result_out[3] ;
wire \alu_result_out[4] ;
wire \alu_result_out[5] ;
wire \alu_result_out[6] ;
wire \alu_result_out[7] ;
wire \alu_result_out[8] ;
wire \alu_result_out[9] ;
wire \alu_result_out[10] ;
wire \alu_result_out[11] ;
wire \alu_result_out[12] ;
wire \alu_result_out[13] ;
wire \alu_result_out[14] ;
wire \alu_result_out[15] ;
wire \alu_result_out[16] ;
wire \alu_result_out[17] ;
wire \alu_result_out[18] ;
wire \alu_result_out[19] ;
wire \alu_result_out[20] ;
wire \alu_result_out[21] ;
wire \alu_result_out[22] ;
wire \alu_result_out[23] ;
wire \alu_result_out[24] ;
wire \alu_result_out[25] ;
wire \alu_result_out[26] ;
wire \alu_result_out[27] ;
wire \alu_result_out[28] ;
wire \alu_result_out[29] ;
wire \alu_result_out[30] ;
wire \alu_result_out[31] ;
wire \ifu_rdata[0] ;
wire \ifu_rdata[1] ;
wire \ifu_rdata[2] ;
wire \ifu_rdata[3] ;
wire \ifu_rdata[4] ;
wire \ifu_rdata[5] ;
wire \ifu_rdata[6] ;
wire \ifu_rdata[7] ;
wire \ifu_rdata[8] ;
wire \ifu_rdata[9] ;
wire \ifu_rdata[10] ;
wire \ifu_rdata[11] ;
wire \ifu_rdata[12] ;
wire \ifu_rdata[13] ;
wire \ifu_rdata[14] ;
wire \ifu_rdata[15] ;
wire \ifu_rdata[16] ;
wire \ifu_rdata[17] ;
wire \ifu_rdata[18] ;
wire \ifu_rdata[19] ;
wire \ifu_rdata[20] ;
wire \ifu_rdata[21] ;
wire \load_data_out[0] ;
wire \load_data_out[1] ;
wire \load_data_out[2] ;
wire \load_data_out[3] ;
wire \load_data_out[4] ;
wire \load_data_out[5] ;
wire \load_data_out[6] ;
wire \load_data_out[7] ;
wire \load_data_out[8] ;
wire \load_data_out[9] ;
wire \load_data_out[10] ;
wire \load_data_out[11] ;
wire \load_data_out[12] ;
wire \load_data_out[13] ;
wire \load_data_out[14] ;
wire \load_data_out[15] ;
wire \load_data_out[16] ;
wire \load_data_out[17] ;
wire \load_data_out[18] ;
wire \load_data_out[19] ;
wire \load_data_out[20] ;
wire \load_data_out[21] ;
wire \load_data_out[22] ;
wire \load_data_out[23] ;
wire \load_data_out[24] ;
wire \load_data_out[25] ;
wire \load_data_out[26] ;
wire \load_data_out[27] ;
wire \load_data_out[28] ;
wire \load_data_out[29] ;
wire \load_data_out[30] ;
wire \load_data_out[31] ;
wire \pc_out[0] ;
wire \pc_out[1] ;
wire \pc_out[2] ;
wire \pc_out[3] ;
wire \pc_out[4] ;
wire \pc_out[5] ;
wire \pc_out[6] ;
wire \pc_out[7] ;
wire \pc_out[8] ;
wire \pc_out[9] ;
wire \pc_out[10] ;
wire \pc_out[11] ;
wire \pc_out[12] ;
wire \pc_out[13] ;
wire \pc_out[14] ;
wire \pc_out[15] ;
wire \pc_out[16] ;
wire \pc_out[17] ;
wire \pc_out[18] ;
wire \pc_out[19] ;
wire \pc_out[20] ;
wire \pc_out[21] ;
wire \pc_out[22] ;
wire \pc_out[23] ;
wire \pc_out[24] ;
wire \pc_out[25] ;
wire \pc_out[26] ;
wire \pc_out[27] ;
wire \pc_out[28] ;
wire \pc_out[29] ;
wire \pc_out[30] ;
wire \pc_out[31] ;
wire \u_lsu.pmem[0] ;
wire \u_lsu.pmem[1] ;
wire \u_lsu.pmem[2] ;
wire \u_lsu.pmem[3] ;
wire \u_lsu.pmem[4] ;
wire \u_lsu.pmem[5] ;
wire \u_lsu.pmem[6] ;
wire \u_lsu.pmem[7] ;
wire \u_lsu.pmem[8] ;
wire \u_lsu.pmem[9] ;
wire \u_lsu.pmem[10] ;
wire \u_lsu.pmem[11] ;
wire \u_lsu.pmem[12] ;
wire \u_lsu.pmem[13] ;
wire \u_lsu.pmem[14] ;
wire \u_lsu.pmem[15] ;
wire \u_lsu.pmem[16] ;
wire \u_lsu.pmem[17] ;
wire \u_lsu.pmem[18] ;
wire \u_lsu.pmem[19] ;
wire \u_lsu.pmem[20] ;
wire \u_lsu.pmem[21] ;
wire \u_lsu.pmem[22] ;
wire \u_lsu.pmem[23] ;
wire \u_lsu.pmem[24] ;
wire \u_lsu.pmem[25] ;
wire \u_lsu.pmem[26] ;
wire \u_lsu.pmem[27] ;
wire \u_lsu.pmem[28] ;
wire \u_lsu.pmem[29] ;
wire \u_lsu.pmem[30] ;
wire \u_lsu.pmem[31] ;
wire \u_lsu.pmem[32] ;
wire \u_lsu.pmem[33] ;
wire \u_lsu.pmem[34] ;
wire \u_lsu.pmem[35] ;
wire \u_lsu.pmem[36] ;
wire \u_lsu.pmem[37] ;
wire \u_lsu.pmem[38] ;
wire \u_lsu.pmem[39] ;
wire \u_lsu.pmem[40] ;
wire \u_lsu.pmem[41] ;
wire \u_lsu.pmem[42] ;
wire \u_lsu.pmem[43] ;
wire \u_lsu.pmem[44] ;
wire \u_lsu.pmem[45] ;
wire \u_lsu.pmem[46] ;
wire \u_lsu.pmem[47] ;
wire \u_lsu.pmem[48] ;
wire \u_lsu.pmem[49] ;
wire \u_lsu.pmem[50] ;
wire \u_lsu.pmem[51] ;
wire \u_lsu.pmem[52] ;
wire \u_lsu.pmem[53] ;
wire \u_lsu.pmem[54] ;
wire \u_lsu.pmem[55] ;
wire \u_lsu.pmem[56] ;
wire \u_lsu.pmem[57] ;
wire \u_lsu.pmem[58] ;
wire \u_lsu.pmem[59] ;
wire \u_lsu.pmem[60] ;
wire \u_lsu.pmem[61] ;
wire \u_lsu.pmem[62] ;
wire \u_lsu.pmem[63] ;
wire \u_lsu.pmem[64] ;
wire \u_lsu.pmem[65] ;
wire \u_lsu.pmem[66] ;
wire \u_lsu.pmem[67] ;
wire \u_lsu.pmem[68] ;
wire \u_lsu.pmem[69] ;
wire \u_lsu.pmem[70] ;
wire \u_lsu.pmem[71] ;
wire \u_lsu.pmem[72] ;
wire \u_lsu.pmem[73] ;
wire \u_lsu.pmem[74] ;
wire \u_lsu.pmem[75] ;
wire \u_lsu.pmem[76] ;
wire \u_lsu.pmem[77] ;
wire \u_lsu.pmem[78] ;
wire \u_lsu.pmem[79] ;
wire \u_lsu.pmem[80] ;
wire \u_lsu.pmem[81] ;
wire \u_lsu.pmem[82] ;
wire \u_lsu.pmem[83] ;
wire \u_lsu.pmem[84] ;
wire \u_lsu.pmem[85] ;
wire \u_lsu.pmem[86] ;
wire \u_lsu.pmem[87] ;
wire \u_lsu.pmem[88] ;
wire \u_lsu.pmem[89] ;
wire \u_lsu.pmem[90] ;
wire \u_lsu.pmem[91] ;
wire \u_lsu.pmem[92] ;
wire \u_lsu.pmem[93] ;
wire \u_lsu.pmem[94] ;
wire \u_lsu.pmem[95] ;
wire \u_lsu.pmem[96] ;
wire \u_lsu.pmem[97] ;
wire \u_lsu.pmem[98] ;
wire \u_lsu.pmem[99] ;
wire \u_lsu.pmem[100] ;
wire \u_lsu.pmem[101] ;
wire \u_lsu.pmem[102] ;
wire \u_lsu.pmem[103] ;
wire \u_lsu.pmem[104] ;
wire \u_lsu.pmem[105] ;
wire \u_lsu.pmem[106] ;
wire \u_lsu.pmem[107] ;
wire \u_lsu.pmem[108] ;
wire \u_lsu.pmem[109] ;
wire \u_lsu.pmem[110] ;
wire \u_lsu.pmem[111] ;
wire \u_lsu.pmem[112] ;
wire \u_lsu.pmem[113] ;
wire \u_lsu.pmem[114] ;
wire \u_lsu.pmem[115] ;
wire \u_lsu.pmem[116] ;
wire \u_lsu.pmem[117] ;
wire \u_lsu.pmem[118] ;
wire \u_lsu.pmem[119] ;
wire \u_lsu.pmem[120] ;
wire \u_lsu.pmem[121] ;
wire \u_lsu.pmem[122] ;
wire \u_lsu.pmem[123] ;
wire \u_lsu.pmem[124] ;
wire \u_lsu.pmem[125] ;
wire \u_lsu.pmem[126] ;
wire \u_lsu.pmem[127] ;
wire \u_lsu.pmem[128] ;
wire \u_lsu.pmem[129] ;
wire \u_lsu.pmem[130] ;
wire \u_lsu.pmem[131] ;
wire \u_lsu.pmem[132] ;
wire \u_lsu.pmem[133] ;
wire \u_lsu.pmem[134] ;
wire \u_lsu.pmem[135] ;
wire \u_lsu.pmem[136] ;
wire \u_lsu.pmem[137] ;
wire \u_lsu.pmem[138] ;
wire \u_lsu.pmem[139] ;
wire \u_lsu.pmem[140] ;
wire \u_lsu.pmem[141] ;
wire \u_lsu.pmem[142] ;
wire \u_lsu.pmem[143] ;
wire \u_lsu.pmem[144] ;
wire \u_lsu.pmem[145] ;
wire \u_lsu.pmem[146] ;
wire \u_lsu.pmem[147] ;
wire \u_lsu.pmem[148] ;
wire \u_lsu.pmem[149] ;
wire \u_lsu.pmem[150] ;
wire \u_lsu.pmem[151] ;
wire \u_lsu.pmem[152] ;
wire \u_lsu.pmem[153] ;
wire \u_lsu.pmem[154] ;
wire \u_lsu.pmem[155] ;
wire \u_lsu.pmem[156] ;
wire \u_lsu.pmem[157] ;
wire \u_lsu.pmem[158] ;
wire \u_lsu.pmem[159] ;
wire \u_lsu.pmem[160] ;
wire \u_lsu.pmem[161] ;
wire \u_lsu.pmem[162] ;
wire \u_lsu.pmem[163] ;
wire \u_lsu.pmem[164] ;
wire \u_lsu.pmem[165] ;
wire \u_lsu.pmem[166] ;
wire \u_lsu.pmem[167] ;
wire \u_lsu.pmem[168] ;
wire \u_lsu.pmem[169] ;
wire \u_lsu.pmem[170] ;
wire \u_lsu.pmem[171] ;
wire \u_lsu.pmem[172] ;
wire \u_lsu.pmem[173] ;
wire \u_lsu.pmem[174] ;
wire \u_lsu.pmem[175] ;
wire \u_lsu.pmem[176] ;
wire \u_lsu.pmem[177] ;
wire \u_lsu.pmem[178] ;
wire \u_lsu.pmem[179] ;
wire \u_lsu.pmem[180] ;
wire \u_lsu.pmem[181] ;
wire \u_lsu.pmem[182] ;
wire \u_lsu.pmem[183] ;
wire \u_lsu.pmem[184] ;
wire \u_lsu.pmem[185] ;
wire \u_lsu.pmem[186] ;
wire \u_lsu.pmem[187] ;
wire \u_lsu.pmem[188] ;
wire \u_lsu.pmem[189] ;
wire \u_lsu.pmem[190] ;
wire \u_lsu.pmem[191] ;
wire \u_lsu.pmem[192] ;
wire \u_lsu.pmem[193] ;
wire \u_lsu.pmem[194] ;
wire \u_lsu.pmem[195] ;
wire \u_lsu.pmem[196] ;
wire \u_lsu.pmem[197] ;
wire \u_lsu.pmem[198] ;
wire \u_lsu.pmem[199] ;
wire \u_lsu.pmem[200] ;
wire \u_lsu.pmem[201] ;
wire \u_lsu.pmem[202] ;
wire \u_lsu.pmem[203] ;
wire \u_lsu.pmem[204] ;
wire \u_lsu.pmem[205] ;
wire \u_lsu.pmem[206] ;
wire \u_lsu.pmem[207] ;
wire \u_lsu.pmem[208] ;
wire \u_lsu.pmem[209] ;
wire \u_lsu.pmem[210] ;
wire \u_lsu.pmem[211] ;
wire \u_lsu.pmem[212] ;
wire \u_lsu.pmem[213] ;
wire \u_lsu.pmem[214] ;
wire \u_lsu.pmem[215] ;
wire \u_lsu.pmem[216] ;
wire \u_lsu.pmem[217] ;
wire \u_lsu.pmem[218] ;
wire \u_lsu.pmem[219] ;
wire \u_lsu.pmem[220] ;
wire \u_lsu.pmem[221] ;
wire \u_lsu.pmem[222] ;
wire \u_lsu.pmem[223] ;
wire \u_lsu.pmem[224] ;
wire \u_lsu.pmem[225] ;
wire \u_lsu.pmem[226] ;
wire \u_lsu.pmem[227] ;
wire \u_lsu.pmem[228] ;
wire \u_lsu.pmem[229] ;
wire \u_lsu.pmem[230] ;
wire \u_lsu.pmem[231] ;
wire \u_lsu.pmem[232] ;
wire \u_lsu.pmem[233] ;
wire \u_lsu.pmem[234] ;
wire \u_lsu.pmem[235] ;
wire \u_lsu.pmem[236] ;
wire \u_lsu.pmem[237] ;
wire \u_lsu.pmem[238] ;
wire \u_lsu.pmem[239] ;
wire \u_lsu.pmem[240] ;
wire \u_lsu.pmem[241] ;
wire \u_lsu.pmem[242] ;
wire \u_lsu.pmem[243] ;
wire \u_lsu.pmem[244] ;
wire \u_lsu.pmem[245] ;
wire \u_lsu.pmem[246] ;
wire \u_lsu.pmem[247] ;
wire \u_lsu.pmem[248] ;
wire \u_lsu.pmem[249] ;
wire \u_lsu.pmem[250] ;
wire \u_lsu.pmem[251] ;
wire \u_lsu.pmem[252] ;
wire \u_lsu.pmem[253] ;
wire \u_lsu.pmem[254] ;
wire \u_lsu.pmem[255] ;
wire \u_lsu.pmem[256] ;
wire \u_lsu.pmem[257] ;
wire \u_lsu.pmem[258] ;
wire \u_lsu.pmem[259] ;
wire \u_lsu.pmem[260] ;
wire \u_lsu.pmem[261] ;
wire \u_lsu.pmem[262] ;
wire \u_lsu.pmem[263] ;
wire \u_lsu.pmem[264] ;
wire \u_lsu.pmem[265] ;
wire \u_lsu.pmem[266] ;
wire \u_lsu.pmem[267] ;
wire \u_lsu.pmem[268] ;
wire \u_lsu.pmem[269] ;
wire \u_lsu.pmem[270] ;
wire \u_lsu.pmem[271] ;
wire \u_lsu.pmem[272] ;
wire \u_lsu.pmem[273] ;
wire \u_lsu.pmem[274] ;
wire \u_lsu.pmem[275] ;
wire \u_lsu.pmem[276] ;
wire \u_lsu.pmem[277] ;
wire \u_lsu.pmem[278] ;
wire \u_lsu.pmem[279] ;
wire \u_lsu.pmem[280] ;
wire \u_lsu.pmem[281] ;
wire \u_lsu.pmem[282] ;
wire \u_lsu.pmem[283] ;
wire \u_lsu.pmem[284] ;
wire \u_lsu.pmem[285] ;
wire \u_lsu.pmem[286] ;
wire \u_lsu.pmem[287] ;
wire \u_lsu.pmem[288] ;
wire \u_lsu.pmem[289] ;
wire \u_lsu.pmem[290] ;
wire \u_lsu.pmem[291] ;
wire \u_lsu.pmem[292] ;
wire \u_lsu.pmem[293] ;
wire \u_lsu.pmem[294] ;
wire \u_lsu.pmem[295] ;
wire \u_lsu.pmem[296] ;
wire \u_lsu.pmem[297] ;
wire \u_lsu.pmem[298] ;
wire \u_lsu.pmem[299] ;
wire \u_lsu.pmem[300] ;
wire \u_lsu.pmem[301] ;
wire \u_lsu.pmem[302] ;
wire \u_lsu.pmem[303] ;
wire \u_lsu.pmem[304] ;
wire \u_lsu.pmem[305] ;
wire \u_lsu.pmem[306] ;
wire \u_lsu.pmem[307] ;
wire \u_lsu.pmem[308] ;
wire \u_lsu.pmem[309] ;
wire \u_lsu.pmem[310] ;
wire \u_lsu.pmem[311] ;
wire \u_lsu.pmem[312] ;
wire \u_lsu.pmem[313] ;
wire \u_lsu.pmem[314] ;
wire \u_lsu.pmem[315] ;
wire \u_lsu.pmem[316] ;
wire \u_lsu.pmem[317] ;
wire \u_lsu.pmem[318] ;
wire \u_lsu.pmem[319] ;
wire \u_lsu.pmem[320] ;
wire \u_lsu.pmem[321] ;
wire \u_lsu.pmem[322] ;
wire \u_lsu.pmem[323] ;
wire \u_lsu.pmem[324] ;
wire \u_lsu.pmem[325] ;
wire \u_lsu.pmem[326] ;
wire \u_lsu.pmem[327] ;
wire \u_lsu.pmem[328] ;
wire \u_lsu.pmem[329] ;
wire \u_lsu.pmem[330] ;
wire \u_lsu.pmem[331] ;
wire \u_lsu.pmem[332] ;
wire \u_lsu.pmem[333] ;
wire \u_lsu.pmem[334] ;
wire \u_lsu.pmem[335] ;
wire \u_lsu.pmem[336] ;
wire \u_lsu.pmem[337] ;
wire \u_lsu.pmem[338] ;
wire \u_lsu.pmem[339] ;
wire \u_lsu.pmem[340] ;
wire \u_lsu.pmem[341] ;
wire \u_lsu.pmem[342] ;
wire \u_lsu.pmem[343] ;
wire \u_lsu.pmem[344] ;
wire \u_lsu.pmem[345] ;
wire \u_lsu.pmem[346] ;
wire \u_lsu.pmem[347] ;
wire \u_lsu.pmem[348] ;
wire \u_lsu.pmem[349] ;
wire \u_lsu.pmem[350] ;
wire \u_lsu.pmem[351] ;
wire \u_lsu.pmem[352] ;
wire \u_lsu.pmem[353] ;
wire \u_lsu.pmem[354] ;
wire \u_lsu.pmem[355] ;
wire \u_lsu.pmem[356] ;
wire \u_lsu.pmem[357] ;
wire \u_lsu.pmem[358] ;
wire \u_lsu.pmem[359] ;
wire \u_lsu.pmem[360] ;
wire \u_lsu.pmem[361] ;
wire \u_lsu.pmem[362] ;
wire \u_lsu.pmem[363] ;
wire \u_lsu.pmem[364] ;
wire \u_lsu.pmem[365] ;
wire \u_lsu.pmem[366] ;
wire \u_lsu.pmem[367] ;
wire \u_lsu.pmem[368] ;
wire \u_lsu.pmem[369] ;
wire \u_lsu.pmem[370] ;
wire \u_lsu.pmem[371] ;
wire \u_lsu.pmem[372] ;
wire \u_lsu.pmem[373] ;
wire \u_lsu.pmem[374] ;
wire \u_lsu.pmem[375] ;
wire \u_lsu.pmem[376] ;
wire \u_lsu.pmem[377] ;
wire \u_lsu.pmem[378] ;
wire \u_lsu.pmem[379] ;
wire \u_lsu.pmem[380] ;
wire \u_lsu.pmem[381] ;
wire \u_lsu.pmem[382] ;
wire \u_lsu.pmem[383] ;
wire \u_lsu.pmem[384] ;
wire \u_lsu.pmem[385] ;
wire \u_lsu.pmem[386] ;
wire \u_lsu.pmem[387] ;
wire \u_lsu.pmem[388] ;
wire \u_lsu.pmem[389] ;
wire \u_lsu.pmem[390] ;
wire \u_lsu.pmem[391] ;
wire \u_lsu.pmem[392] ;
wire \u_lsu.pmem[393] ;
wire \u_lsu.pmem[394] ;
wire \u_lsu.pmem[395] ;
wire \u_lsu.pmem[396] ;
wire \u_lsu.pmem[397] ;
wire \u_lsu.pmem[398] ;
wire \u_lsu.pmem[399] ;
wire \u_lsu.pmem[400] ;
wire \u_lsu.pmem[401] ;
wire \u_lsu.pmem[402] ;
wire \u_lsu.pmem[403] ;
wire \u_lsu.pmem[404] ;
wire \u_lsu.pmem[405] ;
wire \u_lsu.pmem[406] ;
wire \u_lsu.pmem[407] ;
wire \u_lsu.pmem[408] ;
wire \u_lsu.pmem[409] ;
wire \u_lsu.pmem[410] ;
wire \u_lsu.pmem[411] ;
wire \u_lsu.pmem[412] ;
wire \u_lsu.pmem[413] ;
wire \u_lsu.pmem[414] ;
wire \u_lsu.pmem[415] ;
wire \u_lsu.pmem[416] ;
wire \u_lsu.pmem[417] ;
wire \u_lsu.pmem[418] ;
wire \u_lsu.pmem[419] ;
wire \u_lsu.pmem[420] ;
wire \u_lsu.pmem[421] ;
wire \u_lsu.pmem[422] ;
wire \u_lsu.pmem[423] ;
wire \u_lsu.pmem[424] ;
wire \u_lsu.pmem[425] ;
wire \u_lsu.pmem[426] ;
wire \u_lsu.pmem[427] ;
wire \u_lsu.pmem[428] ;
wire \u_lsu.pmem[429] ;
wire \u_lsu.pmem[430] ;
wire \u_lsu.pmem[431] ;
wire \u_lsu.pmem[432] ;
wire \u_lsu.pmem[433] ;
wire \u_lsu.pmem[434] ;
wire \u_lsu.pmem[435] ;
wire \u_lsu.pmem[436] ;
wire \u_lsu.pmem[437] ;
wire \u_lsu.pmem[438] ;
wire \u_lsu.pmem[439] ;
wire \u_lsu.pmem[440] ;
wire \u_lsu.pmem[441] ;
wire \u_lsu.pmem[442] ;
wire \u_lsu.pmem[443] ;
wire \u_lsu.pmem[444] ;
wire \u_lsu.pmem[445] ;
wire \u_lsu.pmem[446] ;
wire \u_lsu.pmem[447] ;
wire \u_lsu.pmem[448] ;
wire \u_lsu.pmem[449] ;
wire \u_lsu.pmem[450] ;
wire \u_lsu.pmem[451] ;
wire \u_lsu.pmem[452] ;
wire \u_lsu.pmem[453] ;
wire \u_lsu.pmem[454] ;
wire \u_lsu.pmem[455] ;
wire \u_lsu.pmem[456] ;
wire \u_lsu.pmem[457] ;
wire \u_lsu.pmem[458] ;
wire \u_lsu.pmem[459] ;
wire \u_lsu.pmem[460] ;
wire \u_lsu.pmem[461] ;
wire \u_lsu.pmem[462] ;
wire \u_lsu.pmem[463] ;
wire \u_lsu.pmem[464] ;
wire \u_lsu.pmem[465] ;
wire \u_lsu.pmem[466] ;
wire \u_lsu.pmem[467] ;
wire \u_lsu.pmem[468] ;
wire \u_lsu.pmem[469] ;
wire \u_lsu.pmem[470] ;
wire \u_lsu.pmem[471] ;
wire \u_lsu.pmem[472] ;
wire \u_lsu.pmem[473] ;
wire \u_lsu.pmem[474] ;
wire \u_lsu.pmem[475] ;
wire \u_lsu.pmem[476] ;
wire \u_lsu.pmem[477] ;
wire \u_lsu.pmem[478] ;
wire \u_lsu.pmem[479] ;
wire \u_lsu.pmem[480] ;
wire \u_lsu.pmem[481] ;
wire \u_lsu.pmem[482] ;
wire \u_lsu.pmem[483] ;
wire \u_lsu.pmem[484] ;
wire \u_lsu.pmem[485] ;
wire \u_lsu.pmem[486] ;
wire \u_lsu.pmem[487] ;
wire \u_lsu.pmem[488] ;
wire \u_lsu.pmem[489] ;
wire \u_lsu.pmem[490] ;
wire \u_lsu.pmem[491] ;
wire \u_lsu.pmem[492] ;
wire \u_lsu.pmem[493] ;
wire \u_lsu.pmem[494] ;
wire \u_lsu.pmem[495] ;
wire \u_lsu.pmem[496] ;
wire \u_lsu.pmem[497] ;
wire \u_lsu.pmem[498] ;
wire \u_lsu.pmem[499] ;
wire \u_lsu.pmem[500] ;
wire \u_lsu.pmem[501] ;
wire \u_lsu.pmem[502] ;
wire \u_lsu.pmem[503] ;
wire \u_lsu.pmem[504] ;
wire \u_lsu.pmem[505] ;
wire \u_lsu.pmem[506] ;
wire \u_lsu.pmem[507] ;
wire \u_lsu.pmem[508] ;
wire \u_lsu.pmem[509] ;
wire \u_lsu.pmem[510] ;
wire \u_lsu.pmem[511] ;
wire \u_lsu.pmem[512] ;
wire \u_lsu.pmem[513] ;
wire \u_lsu.pmem[514] ;
wire \u_lsu.pmem[515] ;
wire \u_lsu.pmem[516] ;
wire \u_lsu.pmem[517] ;
wire \u_lsu.pmem[518] ;
wire \u_lsu.pmem[519] ;
wire \u_lsu.pmem[520] ;
wire \u_lsu.pmem[521] ;
wire \u_lsu.pmem[522] ;
wire \u_lsu.pmem[523] ;
wire \u_lsu.pmem[524] ;
wire \u_lsu.pmem[525] ;
wire \u_lsu.pmem[526] ;
wire \u_lsu.pmem[527] ;
wire \u_lsu.pmem[528] ;
wire \u_lsu.pmem[529] ;
wire \u_lsu.pmem[530] ;
wire \u_lsu.pmem[531] ;
wire \u_lsu.pmem[532] ;
wire \u_lsu.pmem[533] ;
wire \u_lsu.pmem[534] ;
wire \u_lsu.pmem[535] ;
wire \u_lsu.pmem[536] ;
wire \u_lsu.pmem[537] ;
wire \u_lsu.pmem[538] ;
wire \u_lsu.pmem[539] ;
wire \u_lsu.pmem[540] ;
wire \u_lsu.pmem[541] ;
wire \u_lsu.pmem[542] ;
wire \u_lsu.pmem[543] ;
wire \u_lsu.pmem[544] ;
wire \u_lsu.pmem[545] ;
wire \u_lsu.pmem[546] ;
wire \u_lsu.pmem[547] ;
wire \u_lsu.pmem[548] ;
wire \u_lsu.pmem[549] ;
wire \u_lsu.pmem[550] ;
wire \u_lsu.pmem[551] ;
wire \u_lsu.pmem[552] ;
wire \u_lsu.pmem[553] ;
wire \u_lsu.pmem[554] ;
wire \u_lsu.pmem[555] ;
wire \u_lsu.pmem[556] ;
wire \u_lsu.pmem[557] ;
wire \u_lsu.pmem[558] ;
wire \u_lsu.pmem[559] ;
wire \u_lsu.pmem[560] ;
wire \u_lsu.pmem[561] ;
wire \u_lsu.pmem[562] ;
wire \u_lsu.pmem[563] ;
wire \u_lsu.pmem[564] ;
wire \u_lsu.pmem[565] ;
wire \u_lsu.pmem[566] ;
wire \u_lsu.pmem[567] ;
wire \u_lsu.pmem[568] ;
wire \u_lsu.pmem[569] ;
wire \u_lsu.pmem[570] ;
wire \u_lsu.pmem[571] ;
wire \u_lsu.pmem[572] ;
wire \u_lsu.pmem[573] ;
wire \u_lsu.pmem[574] ;
wire \u_lsu.pmem[575] ;
wire \u_lsu.pmem[576] ;
wire \u_lsu.pmem[577] ;
wire \u_lsu.pmem[578] ;
wire \u_lsu.pmem[579] ;
wire \u_lsu.pmem[580] ;
wire \u_lsu.pmem[581] ;
wire \u_lsu.pmem[582] ;
wire \u_lsu.pmem[583] ;
wire \u_lsu.pmem[584] ;
wire \u_lsu.pmem[585] ;
wire \u_lsu.pmem[586] ;
wire \u_lsu.pmem[587] ;
wire \u_lsu.pmem[588] ;
wire \u_lsu.pmem[589] ;
wire \u_lsu.pmem[590] ;
wire \u_lsu.pmem[591] ;
wire \u_lsu.pmem[592] ;
wire \u_lsu.pmem[593] ;
wire \u_lsu.pmem[594] ;
wire \u_lsu.pmem[595] ;
wire \u_lsu.pmem[596] ;
wire \u_lsu.pmem[597] ;
wire \u_lsu.pmem[598] ;
wire \u_lsu.pmem[599] ;
wire \u_lsu.pmem[600] ;
wire \u_lsu.pmem[601] ;
wire \u_lsu.pmem[602] ;
wire \u_lsu.pmem[603] ;
wire \u_lsu.pmem[604] ;
wire \u_lsu.pmem[605] ;
wire \u_lsu.pmem[606] ;
wire \u_lsu.pmem[607] ;
wire \u_lsu.pmem[608] ;
wire \u_lsu.pmem[609] ;
wire \u_lsu.pmem[610] ;
wire \u_lsu.pmem[611] ;
wire \u_lsu.pmem[612] ;
wire \u_lsu.pmem[613] ;
wire \u_lsu.pmem[614] ;
wire \u_lsu.pmem[615] ;
wire \u_lsu.pmem[616] ;
wire \u_lsu.pmem[617] ;
wire \u_lsu.pmem[618] ;
wire \u_lsu.pmem[619] ;
wire \u_lsu.pmem[620] ;
wire \u_lsu.pmem[621] ;
wire \u_lsu.pmem[622] ;
wire \u_lsu.pmem[623] ;
wire \u_lsu.pmem[624] ;
wire \u_lsu.pmem[625] ;
wire \u_lsu.pmem[626] ;
wire \u_lsu.pmem[627] ;
wire \u_lsu.pmem[628] ;
wire \u_lsu.pmem[629] ;
wire \u_lsu.pmem[630] ;
wire \u_lsu.pmem[631] ;
wire \u_lsu.pmem[632] ;
wire \u_lsu.pmem[633] ;
wire \u_lsu.pmem[634] ;
wire \u_lsu.pmem[635] ;
wire \u_lsu.pmem[636] ;
wire \u_lsu.pmem[637] ;
wire \u_lsu.pmem[638] ;
wire \u_lsu.pmem[639] ;
wire \u_lsu.pmem[640] ;
wire \u_lsu.pmem[641] ;
wire \u_lsu.pmem[642] ;
wire \u_lsu.pmem[643] ;
wire \u_lsu.pmem[644] ;
wire \u_lsu.pmem[645] ;
wire \u_lsu.pmem[646] ;
wire \u_lsu.pmem[647] ;
wire \u_lsu.pmem[648] ;
wire \u_lsu.pmem[649] ;
wire \u_lsu.pmem[650] ;
wire \u_lsu.pmem[651] ;
wire \u_lsu.pmem[652] ;
wire \u_lsu.pmem[653] ;
wire \u_lsu.pmem[654] ;
wire \u_lsu.pmem[655] ;
wire \u_lsu.pmem[656] ;
wire \u_lsu.pmem[657] ;
wire \u_lsu.pmem[658] ;
wire \u_lsu.pmem[659] ;
wire \u_lsu.pmem[660] ;
wire \u_lsu.pmem[661] ;
wire \u_lsu.pmem[662] ;
wire \u_lsu.pmem[663] ;
wire \u_lsu.pmem[664] ;
wire \u_lsu.pmem[665] ;
wire \u_lsu.pmem[666] ;
wire \u_lsu.pmem[667] ;
wire \u_lsu.pmem[668] ;
wire \u_lsu.pmem[669] ;
wire \u_lsu.pmem[670] ;
wire \u_lsu.pmem[671] ;
wire \u_lsu.pmem[672] ;
wire \u_lsu.pmem[673] ;
wire \u_lsu.pmem[674] ;
wire \u_lsu.pmem[675] ;
wire \u_lsu.pmem[676] ;
wire \u_lsu.pmem[677] ;
wire \u_lsu.pmem[678] ;
wire \u_lsu.pmem[679] ;
wire \u_lsu.pmem[680] ;
wire \u_lsu.pmem[681] ;
wire \u_lsu.pmem[682] ;
wire \u_lsu.pmem[683] ;
wire \u_lsu.pmem[684] ;
wire \u_lsu.pmem[685] ;
wire \u_lsu.pmem[686] ;
wire \u_lsu.pmem[687] ;
wire \u_lsu.pmem[688] ;
wire \u_lsu.pmem[689] ;
wire \u_lsu.pmem[690] ;
wire \u_lsu.pmem[691] ;
wire \u_lsu.pmem[692] ;
wire \u_lsu.pmem[693] ;
wire \u_lsu.pmem[694] ;
wire \u_lsu.pmem[695] ;
wire \u_lsu.pmem[696] ;
wire \u_lsu.pmem[697] ;
wire \u_lsu.pmem[698] ;
wire \u_lsu.pmem[699] ;
wire \u_lsu.pmem[700] ;
wire \u_lsu.pmem[701] ;
wire \u_lsu.pmem[702] ;
wire \u_lsu.pmem[703] ;
wire \u_lsu.pmem[704] ;
wire \u_lsu.pmem[705] ;
wire \u_lsu.pmem[706] ;
wire \u_lsu.pmem[707] ;
wire \u_lsu.pmem[708] ;
wire \u_lsu.pmem[709] ;
wire \u_lsu.pmem[710] ;
wire \u_lsu.pmem[711] ;
wire \u_lsu.pmem[712] ;
wire \u_lsu.pmem[713] ;
wire \u_lsu.pmem[714] ;
wire \u_lsu.pmem[715] ;
wire \u_lsu.pmem[716] ;
wire \u_lsu.pmem[717] ;
wire \u_lsu.pmem[718] ;
wire \u_lsu.pmem[719] ;
wire \u_lsu.pmem[720] ;
wire \u_lsu.pmem[721] ;
wire \u_lsu.pmem[722] ;
wire \u_lsu.pmem[723] ;
wire \u_lsu.pmem[724] ;
wire \u_lsu.pmem[725] ;
wire \u_lsu.pmem[726] ;
wire \u_lsu.pmem[727] ;
wire \u_lsu.pmem[728] ;
wire \u_lsu.pmem[729] ;
wire \u_lsu.pmem[730] ;
wire \u_lsu.pmem[731] ;
wire \u_lsu.pmem[732] ;
wire \u_lsu.pmem[733] ;
wire \u_lsu.pmem[734] ;
wire \u_lsu.pmem[735] ;
wire \u_lsu.pmem[736] ;
wire \u_lsu.pmem[737] ;
wire \u_lsu.pmem[738] ;
wire \u_lsu.pmem[739] ;
wire \u_lsu.pmem[740] ;
wire \u_lsu.pmem[741] ;
wire \u_lsu.pmem[742] ;
wire \u_lsu.pmem[743] ;
wire \u_lsu.pmem[744] ;
wire \u_lsu.pmem[745] ;
wire \u_lsu.pmem[746] ;
wire \u_lsu.pmem[747] ;
wire \u_lsu.pmem[748] ;
wire \u_lsu.pmem[749] ;
wire \u_lsu.pmem[750] ;
wire \u_lsu.pmem[751] ;
wire \u_lsu.pmem[752] ;
wire \u_lsu.pmem[753] ;
wire \u_lsu.pmem[754] ;
wire \u_lsu.pmem[755] ;
wire \u_lsu.pmem[756] ;
wire \u_lsu.pmem[757] ;
wire \u_lsu.pmem[758] ;
wire \u_lsu.pmem[759] ;
wire \u_lsu.pmem[760] ;
wire \u_lsu.pmem[761] ;
wire \u_lsu.pmem[762] ;
wire \u_lsu.pmem[763] ;
wire \u_lsu.pmem[764] ;
wire \u_lsu.pmem[765] ;
wire \u_lsu.pmem[766] ;
wire \u_lsu.pmem[767] ;
wire \u_lsu.pmem[768] ;
wire \u_lsu.pmem[769] ;
wire \u_lsu.pmem[770] ;
wire \u_lsu.pmem[771] ;
wire \u_lsu.pmem[772] ;
wire \u_lsu.pmem[773] ;
wire \u_lsu.pmem[774] ;
wire \u_lsu.pmem[775] ;
wire \u_lsu.pmem[776] ;
wire \u_lsu.pmem[777] ;
wire \u_lsu.pmem[778] ;
wire \u_lsu.pmem[779] ;
wire \u_lsu.pmem[780] ;
wire \u_lsu.pmem[781] ;
wire \u_lsu.pmem[782] ;
wire \u_lsu.pmem[783] ;
wire \u_lsu.pmem[784] ;
wire \u_lsu.pmem[785] ;
wire \u_lsu.pmem[786] ;
wire \u_lsu.pmem[787] ;
wire \u_lsu.pmem[788] ;
wire \u_lsu.pmem[789] ;
wire \u_lsu.pmem[790] ;
wire \u_lsu.pmem[791] ;
wire \u_lsu.pmem[792] ;
wire \u_lsu.pmem[793] ;
wire \u_lsu.pmem[794] ;
wire \u_lsu.pmem[795] ;
wire \u_lsu.pmem[796] ;
wire \u_lsu.pmem[797] ;
wire \u_lsu.pmem[798] ;
wire \u_lsu.pmem[799] ;
wire \u_lsu.pmem[800] ;
wire \u_lsu.pmem[801] ;
wire \u_lsu.pmem[802] ;
wire \u_lsu.pmem[803] ;
wire \u_lsu.pmem[804] ;
wire \u_lsu.pmem[805] ;
wire \u_lsu.pmem[806] ;
wire \u_lsu.pmem[807] ;
wire \u_lsu.pmem[808] ;
wire \u_lsu.pmem[809] ;
wire \u_lsu.pmem[810] ;
wire \u_lsu.pmem[811] ;
wire \u_lsu.pmem[812] ;
wire \u_lsu.pmem[813] ;
wire \u_lsu.pmem[814] ;
wire \u_lsu.pmem[815] ;
wire \u_lsu.pmem[816] ;
wire \u_lsu.pmem[817] ;
wire \u_lsu.pmem[818] ;
wire \u_lsu.pmem[819] ;
wire \u_lsu.pmem[820] ;
wire \u_lsu.pmem[821] ;
wire \u_lsu.pmem[822] ;
wire \u_lsu.pmem[823] ;
wire \u_lsu.pmem[824] ;
wire \u_lsu.pmem[825] ;
wire \u_lsu.pmem[826] ;
wire \u_lsu.pmem[827] ;
wire \u_lsu.pmem[828] ;
wire \u_lsu.pmem[829] ;
wire \u_lsu.pmem[830] ;
wire \u_lsu.pmem[831] ;
wire \u_lsu.pmem[832] ;
wire \u_lsu.pmem[833] ;
wire \u_lsu.pmem[834] ;
wire \u_lsu.pmem[835] ;
wire \u_lsu.pmem[836] ;
wire \u_lsu.pmem[837] ;
wire \u_lsu.pmem[838] ;
wire \u_lsu.pmem[839] ;
wire \u_lsu.pmem[840] ;
wire \u_lsu.pmem[841] ;
wire \u_lsu.pmem[842] ;
wire \u_lsu.pmem[843] ;
wire \u_lsu.pmem[844] ;
wire \u_lsu.pmem[845] ;
wire \u_lsu.pmem[846] ;
wire \u_lsu.pmem[847] ;
wire \u_lsu.pmem[848] ;
wire \u_lsu.pmem[849] ;
wire \u_lsu.pmem[850] ;
wire \u_lsu.pmem[851] ;
wire \u_lsu.pmem[852] ;
wire \u_lsu.pmem[853] ;
wire \u_lsu.pmem[854] ;
wire \u_lsu.pmem[855] ;
wire \u_lsu.pmem[856] ;
wire \u_lsu.pmem[857] ;
wire \u_lsu.pmem[858] ;
wire \u_lsu.pmem[859] ;
wire \u_lsu.pmem[860] ;
wire \u_lsu.pmem[861] ;
wire \u_lsu.pmem[862] ;
wire \u_lsu.pmem[863] ;
wire \u_lsu.pmem[864] ;
wire \u_lsu.pmem[865] ;
wire \u_lsu.pmem[866] ;
wire \u_lsu.pmem[867] ;
wire \u_lsu.pmem[868] ;
wire \u_lsu.pmem[869] ;
wire \u_lsu.pmem[870] ;
wire \u_lsu.pmem[871] ;
wire \u_lsu.pmem[872] ;
wire \u_lsu.pmem[873] ;
wire \u_lsu.pmem[874] ;
wire \u_lsu.pmem[875] ;
wire \u_lsu.pmem[876] ;
wire \u_lsu.pmem[877] ;
wire \u_lsu.pmem[878] ;
wire \u_lsu.pmem[879] ;
wire \u_lsu.pmem[880] ;
wire \u_lsu.pmem[881] ;
wire \u_lsu.pmem[882] ;
wire \u_lsu.pmem[883] ;
wire \u_lsu.pmem[884] ;
wire \u_lsu.pmem[885] ;
wire \u_lsu.pmem[886] ;
wire \u_lsu.pmem[887] ;
wire \u_lsu.pmem[888] ;
wire \u_lsu.pmem[889] ;
wire \u_lsu.pmem[890] ;
wire \u_lsu.pmem[891] ;
wire \u_lsu.pmem[892] ;
wire \u_lsu.pmem[893] ;
wire \u_lsu.pmem[894] ;
wire \u_lsu.pmem[895] ;
wire \u_lsu.pmem[896] ;
wire \u_lsu.pmem[897] ;
wire \u_lsu.pmem[898] ;
wire \u_lsu.pmem[899] ;
wire \u_lsu.pmem[900] ;
wire \u_lsu.pmem[901] ;
wire \u_lsu.pmem[902] ;
wire \u_lsu.pmem[903] ;
wire \u_lsu.pmem[904] ;
wire \u_lsu.pmem[905] ;
wire \u_lsu.pmem[906] ;
wire \u_lsu.pmem[907] ;
wire \u_lsu.pmem[908] ;
wire \u_lsu.pmem[909] ;
wire \u_lsu.pmem[910] ;
wire \u_lsu.pmem[911] ;
wire \u_lsu.pmem[912] ;
wire \u_lsu.pmem[913] ;
wire \u_lsu.pmem[914] ;
wire \u_lsu.pmem[915] ;
wire \u_lsu.pmem[916] ;
wire \u_lsu.pmem[917] ;
wire \u_lsu.pmem[918] ;
wire \u_lsu.pmem[919] ;
wire \u_lsu.pmem[920] ;
wire \u_lsu.pmem[921] ;
wire \u_lsu.pmem[922] ;
wire \u_lsu.pmem[923] ;
wire \u_lsu.pmem[924] ;
wire \u_lsu.pmem[925] ;
wire \u_lsu.pmem[926] ;
wire \u_lsu.pmem[927] ;
wire \u_lsu.pmem[928] ;
wire \u_lsu.pmem[929] ;
wire \u_lsu.pmem[930] ;
wire \u_lsu.pmem[931] ;
wire \u_lsu.pmem[932] ;
wire \u_lsu.pmem[933] ;
wire \u_lsu.pmem[934] ;
wire \u_lsu.pmem[935] ;
wire \u_lsu.pmem[936] ;
wire \u_lsu.pmem[937] ;
wire \u_lsu.pmem[938] ;
wire \u_lsu.pmem[939] ;
wire \u_lsu.pmem[940] ;
wire \u_lsu.pmem[941] ;
wire \u_lsu.pmem[942] ;
wire \u_lsu.pmem[943] ;
wire \u_lsu.pmem[944] ;
wire \u_lsu.pmem[945] ;
wire \u_lsu.pmem[946] ;
wire \u_lsu.pmem[947] ;
wire \u_lsu.pmem[948] ;
wire \u_lsu.pmem[949] ;
wire \u_lsu.pmem[950] ;
wire \u_lsu.pmem[951] ;
wire \u_lsu.pmem[952] ;
wire \u_lsu.pmem[953] ;
wire \u_lsu.pmem[954] ;
wire \u_lsu.pmem[955] ;
wire \u_lsu.pmem[956] ;
wire \u_lsu.pmem[957] ;
wire \u_lsu.pmem[958] ;
wire \u_lsu.pmem[959] ;
wire \u_lsu.pmem[960] ;
wire \u_lsu.pmem[961] ;
wire \u_lsu.pmem[962] ;
wire \u_lsu.pmem[963] ;
wire \u_lsu.pmem[964] ;
wire \u_lsu.pmem[965] ;
wire \u_lsu.pmem[966] ;
wire \u_lsu.pmem[967] ;
wire \u_lsu.pmem[968] ;
wire \u_lsu.pmem[969] ;
wire \u_lsu.pmem[970] ;
wire \u_lsu.pmem[971] ;
wire \u_lsu.pmem[972] ;
wire \u_lsu.pmem[973] ;
wire \u_lsu.pmem[974] ;
wire \u_lsu.pmem[975] ;
wire \u_lsu.pmem[976] ;
wire \u_lsu.pmem[977] ;
wire \u_lsu.pmem[978] ;
wire \u_lsu.pmem[979] ;
wire \u_lsu.pmem[980] ;
wire \u_lsu.pmem[981] ;
wire \u_lsu.pmem[982] ;
wire \u_lsu.pmem[983] ;
wire \u_lsu.pmem[984] ;
wire \u_lsu.pmem[985] ;
wire \u_lsu.pmem[986] ;
wire \u_lsu.pmem[987] ;
wire \u_lsu.pmem[988] ;
wire \u_lsu.pmem[989] ;
wire \u_lsu.pmem[990] ;
wire \u_lsu.pmem[991] ;
wire \u_lsu.pmem[992] ;
wire \u_lsu.pmem[993] ;
wire \u_lsu.pmem[994] ;
wire \u_lsu.pmem[995] ;
wire \u_lsu.pmem[996] ;
wire \u_lsu.pmem[997] ;
wire \u_lsu.pmem[998] ;
wire \u_lsu.pmem[999] ;
wire \u_lsu.pmem[1000] ;
wire \u_lsu.pmem[1001] ;
wire \u_lsu.pmem[1002] ;
wire \u_lsu.pmem[1003] ;
wire \u_lsu.pmem[1004] ;
wire \u_lsu.pmem[1005] ;
wire \u_lsu.pmem[1006] ;
wire \u_lsu.pmem[1007] ;
wire \u_lsu.pmem[1008] ;
wire \u_lsu.pmem[1009] ;
wire \u_lsu.pmem[1010] ;
wire \u_lsu.pmem[1011] ;
wire \u_lsu.pmem[1012] ;
wire \u_lsu.pmem[1013] ;
wire \u_lsu.pmem[1014] ;
wire \u_lsu.pmem[1015] ;
wire \u_lsu.pmem[1016] ;
wire \u_lsu.pmem[1017] ;
wire \u_lsu.pmem[1018] ;
wire \u_lsu.pmem[1019] ;
wire \u_lsu.pmem[1020] ;
wire \u_lsu.pmem[1021] ;
wire \u_lsu.pmem[1022] ;
wire \u_lsu.pmem[1023] ;
wire \u_lsu.pmem[1024] ;
wire \u_lsu.pmem[1025] ;
wire \u_lsu.pmem[1026] ;
wire \u_lsu.pmem[1027] ;
wire \u_lsu.pmem[1028] ;
wire \u_lsu.pmem[1029] ;
wire \u_lsu.pmem[1030] ;
wire \u_lsu.pmem[1031] ;
wire \u_lsu.pmem[1032] ;
wire \u_lsu.pmem[1033] ;
wire \u_lsu.pmem[1034] ;
wire \u_lsu.pmem[1035] ;
wire \u_lsu.pmem[1036] ;
wire \u_lsu.pmem[1037] ;
wire \u_lsu.pmem[1038] ;
wire \u_lsu.pmem[1039] ;
wire \u_lsu.pmem[1040] ;
wire \u_lsu.pmem[1041] ;
wire \u_lsu.pmem[1042] ;
wire \u_lsu.pmem[1043] ;
wire \u_lsu.pmem[1044] ;
wire \u_lsu.pmem[1045] ;
wire \u_lsu.pmem[1046] ;
wire \u_lsu.pmem[1047] ;
wire \u_lsu.pmem[1048] ;
wire \u_lsu.pmem[1049] ;
wire \u_lsu.pmem[1050] ;
wire \u_lsu.pmem[1051] ;
wire \u_lsu.pmem[1052] ;
wire \u_lsu.pmem[1053] ;
wire \u_lsu.pmem[1054] ;
wire \u_lsu.pmem[1055] ;
wire \u_lsu.pmem[1056] ;
wire \u_lsu.pmem[1057] ;
wire \u_lsu.pmem[1058] ;
wire \u_lsu.pmem[1059] ;
wire \u_lsu.pmem[1060] ;
wire \u_lsu.pmem[1061] ;
wire \u_lsu.pmem[1062] ;
wire \u_lsu.pmem[1063] ;
wire \u_lsu.pmem[1064] ;
wire \u_lsu.pmem[1065] ;
wire \u_lsu.pmem[1066] ;
wire \u_lsu.pmem[1067] ;
wire \u_lsu.pmem[1068] ;
wire \u_lsu.pmem[1069] ;
wire \u_lsu.pmem[1070] ;
wire \u_lsu.pmem[1071] ;
wire \u_lsu.pmem[1072] ;
wire \u_lsu.pmem[1073] ;
wire \u_lsu.pmem[1074] ;
wire \u_lsu.pmem[1075] ;
wire \u_lsu.pmem[1076] ;
wire \u_lsu.pmem[1077] ;
wire \u_lsu.pmem[1078] ;
wire \u_lsu.pmem[1079] ;
wire \u_lsu.pmem[1080] ;
wire \u_lsu.pmem[1081] ;
wire \u_lsu.pmem[1082] ;
wire \u_lsu.pmem[1083] ;
wire \u_lsu.pmem[1084] ;
wire \u_lsu.pmem[1085] ;
wire \u_lsu.pmem[1086] ;
wire \u_lsu.pmem[1087] ;
wire \u_lsu.pmem[1088] ;
wire \u_lsu.pmem[1089] ;
wire \u_lsu.pmem[1090] ;
wire \u_lsu.pmem[1091] ;
wire \u_lsu.pmem[1092] ;
wire \u_lsu.pmem[1093] ;
wire \u_lsu.pmem[1094] ;
wire \u_lsu.pmem[1095] ;
wire \u_lsu.pmem[1096] ;
wire \u_lsu.pmem[1097] ;
wire \u_lsu.pmem[1098] ;
wire \u_lsu.pmem[1099] ;
wire \u_lsu.pmem[1100] ;
wire \u_lsu.pmem[1101] ;
wire \u_lsu.pmem[1102] ;
wire \u_lsu.pmem[1103] ;
wire \u_lsu.pmem[1104] ;
wire \u_lsu.pmem[1105] ;
wire \u_lsu.pmem[1106] ;
wire \u_lsu.pmem[1107] ;
wire \u_lsu.pmem[1108] ;
wire \u_lsu.pmem[1109] ;
wire \u_lsu.pmem[1110] ;
wire \u_lsu.pmem[1111] ;
wire \u_lsu.pmem[1112] ;
wire \u_lsu.pmem[1113] ;
wire \u_lsu.pmem[1114] ;
wire \u_lsu.pmem[1115] ;
wire \u_lsu.pmem[1116] ;
wire \u_lsu.pmem[1117] ;
wire \u_lsu.pmem[1118] ;
wire \u_lsu.pmem[1119] ;
wire \u_lsu.pmem[1120] ;
wire \u_lsu.pmem[1121] ;
wire \u_lsu.pmem[1122] ;
wire \u_lsu.pmem[1123] ;
wire \u_lsu.pmem[1124] ;
wire \u_lsu.pmem[1125] ;
wire \u_lsu.pmem[1126] ;
wire \u_lsu.pmem[1127] ;
wire \u_lsu.pmem[1128] ;
wire \u_lsu.pmem[1129] ;
wire \u_lsu.pmem[1130] ;
wire \u_lsu.pmem[1131] ;
wire \u_lsu.pmem[1132] ;
wire \u_lsu.pmem[1133] ;
wire \u_lsu.pmem[1134] ;
wire \u_lsu.pmem[1135] ;
wire \u_lsu.pmem[1136] ;
wire \u_lsu.pmem[1137] ;
wire \u_lsu.pmem[1138] ;
wire \u_lsu.pmem[1139] ;
wire \u_lsu.pmem[1140] ;
wire \u_lsu.pmem[1141] ;
wire \u_lsu.pmem[1142] ;
wire \u_lsu.pmem[1143] ;
wire \u_lsu.pmem[1144] ;
wire \u_lsu.pmem[1145] ;
wire \u_lsu.pmem[1146] ;
wire \u_lsu.pmem[1147] ;
wire \u_lsu.pmem[1148] ;
wire \u_lsu.pmem[1149] ;
wire \u_lsu.pmem[1150] ;
wire \u_lsu.pmem[1151] ;
wire \u_lsu.pmem[1152] ;
wire \u_lsu.pmem[1153] ;
wire \u_lsu.pmem[1154] ;
wire \u_lsu.pmem[1155] ;
wire \u_lsu.pmem[1156] ;
wire \u_lsu.pmem[1157] ;
wire \u_lsu.pmem[1158] ;
wire \u_lsu.pmem[1159] ;
wire \u_lsu.pmem[1160] ;
wire \u_lsu.pmem[1161] ;
wire \u_lsu.pmem[1162] ;
wire \u_lsu.pmem[1163] ;
wire \u_lsu.pmem[1164] ;
wire \u_lsu.pmem[1165] ;
wire \u_lsu.pmem[1166] ;
wire \u_lsu.pmem[1167] ;
wire \u_lsu.pmem[1168] ;
wire \u_lsu.pmem[1169] ;
wire \u_lsu.pmem[1170] ;
wire \u_lsu.pmem[1171] ;
wire \u_lsu.pmem[1172] ;
wire \u_lsu.pmem[1173] ;
wire \u_lsu.pmem[1174] ;
wire \u_lsu.pmem[1175] ;
wire \u_lsu.pmem[1176] ;
wire \u_lsu.pmem[1177] ;
wire \u_lsu.pmem[1178] ;
wire \u_lsu.pmem[1179] ;
wire \u_lsu.pmem[1180] ;
wire \u_lsu.pmem[1181] ;
wire \u_lsu.pmem[1182] ;
wire \u_lsu.pmem[1183] ;
wire \u_lsu.pmem[1184] ;
wire \u_lsu.pmem[1185] ;
wire \u_lsu.pmem[1186] ;
wire \u_lsu.pmem[1187] ;
wire \u_lsu.pmem[1188] ;
wire \u_lsu.pmem[1189] ;
wire \u_lsu.pmem[1190] ;
wire \u_lsu.pmem[1191] ;
wire \u_lsu.pmem[1192] ;
wire \u_lsu.pmem[1193] ;
wire \u_lsu.pmem[1194] ;
wire \u_lsu.pmem[1195] ;
wire \u_lsu.pmem[1196] ;
wire \u_lsu.pmem[1197] ;
wire \u_lsu.pmem[1198] ;
wire \u_lsu.pmem[1199] ;
wire \u_lsu.pmem[1200] ;
wire \u_lsu.pmem[1201] ;
wire \u_lsu.pmem[1202] ;
wire \u_lsu.pmem[1203] ;
wire \u_lsu.pmem[1204] ;
wire \u_lsu.pmem[1205] ;
wire \u_lsu.pmem[1206] ;
wire \u_lsu.pmem[1207] ;
wire \u_lsu.pmem[1208] ;
wire \u_lsu.pmem[1209] ;
wire \u_lsu.pmem[1210] ;
wire \u_lsu.pmem[1211] ;
wire \u_lsu.pmem[1212] ;
wire \u_lsu.pmem[1213] ;
wire \u_lsu.pmem[1214] ;
wire \u_lsu.pmem[1215] ;
wire \u_lsu.pmem[1216] ;
wire \u_lsu.pmem[1217] ;
wire \u_lsu.pmem[1218] ;
wire \u_lsu.pmem[1219] ;
wire \u_lsu.pmem[1220] ;
wire \u_lsu.pmem[1221] ;
wire \u_lsu.pmem[1222] ;
wire \u_lsu.pmem[1223] ;
wire \u_lsu.pmem[1224] ;
wire \u_lsu.pmem[1225] ;
wire \u_lsu.pmem[1226] ;
wire \u_lsu.pmem[1227] ;
wire \u_lsu.pmem[1228] ;
wire \u_lsu.pmem[1229] ;
wire \u_lsu.pmem[1230] ;
wire \u_lsu.pmem[1231] ;
wire \u_lsu.pmem[1232] ;
wire \u_lsu.pmem[1233] ;
wire \u_lsu.pmem[1234] ;
wire \u_lsu.pmem[1235] ;
wire \u_lsu.pmem[1236] ;
wire \u_lsu.pmem[1237] ;
wire \u_lsu.pmem[1238] ;
wire \u_lsu.pmem[1239] ;
wire \u_lsu.pmem[1240] ;
wire \u_lsu.pmem[1241] ;
wire \u_lsu.pmem[1242] ;
wire \u_lsu.pmem[1243] ;
wire \u_lsu.pmem[1244] ;
wire \u_lsu.pmem[1245] ;
wire \u_lsu.pmem[1246] ;
wire \u_lsu.pmem[1247] ;
wire \u_lsu.pmem[1248] ;
wire \u_lsu.pmem[1249] ;
wire \u_lsu.pmem[1250] ;
wire \u_lsu.pmem[1251] ;
wire \u_lsu.pmem[1252] ;
wire \u_lsu.pmem[1253] ;
wire \u_lsu.pmem[1254] ;
wire \u_lsu.pmem[1255] ;
wire \u_lsu.pmem[1256] ;
wire \u_lsu.pmem[1257] ;
wire \u_lsu.pmem[1258] ;
wire \u_lsu.pmem[1259] ;
wire \u_lsu.pmem[1260] ;
wire \u_lsu.pmem[1261] ;
wire \u_lsu.pmem[1262] ;
wire \u_lsu.pmem[1263] ;
wire \u_lsu.pmem[1264] ;
wire \u_lsu.pmem[1265] ;
wire \u_lsu.pmem[1266] ;
wire \u_lsu.pmem[1267] ;
wire \u_lsu.pmem[1268] ;
wire \u_lsu.pmem[1269] ;
wire \u_lsu.pmem[1270] ;
wire \u_lsu.pmem[1271] ;
wire \u_lsu.pmem[1272] ;
wire \u_lsu.pmem[1273] ;
wire \u_lsu.pmem[1274] ;
wire \u_lsu.pmem[1275] ;
wire \u_lsu.pmem[1276] ;
wire \u_lsu.pmem[1277] ;
wire \u_lsu.pmem[1278] ;
wire \u_lsu.pmem[1279] ;
wire \u_lsu.pmem[1280] ;
wire \u_lsu.pmem[1281] ;
wire \u_lsu.pmem[1282] ;
wire \u_lsu.pmem[1283] ;
wire \u_lsu.pmem[1284] ;
wire \u_lsu.pmem[1285] ;
wire \u_lsu.pmem[1286] ;
wire \u_lsu.pmem[1287] ;
wire \u_lsu.pmem[1288] ;
wire \u_lsu.pmem[1289] ;
wire \u_lsu.pmem[1290] ;
wire \u_lsu.pmem[1291] ;
wire \u_lsu.pmem[1292] ;
wire \u_lsu.pmem[1293] ;
wire \u_lsu.pmem[1294] ;
wire \u_lsu.pmem[1295] ;
wire \u_lsu.pmem[1296] ;
wire \u_lsu.pmem[1297] ;
wire \u_lsu.pmem[1298] ;
wire \u_lsu.pmem[1299] ;
wire \u_lsu.pmem[1300] ;
wire \u_lsu.pmem[1301] ;
wire \u_lsu.pmem[1302] ;
wire \u_lsu.pmem[1303] ;
wire \u_lsu.pmem[1304] ;
wire \u_lsu.pmem[1305] ;
wire \u_lsu.pmem[1306] ;
wire \u_lsu.pmem[1307] ;
wire \u_lsu.pmem[1308] ;
wire \u_lsu.pmem[1309] ;
wire \u_lsu.pmem[1310] ;
wire \u_lsu.pmem[1311] ;
wire \u_lsu.pmem[1312] ;
wire \u_lsu.pmem[1313] ;
wire \u_lsu.pmem[1314] ;
wire \u_lsu.pmem[1315] ;
wire \u_lsu.pmem[1316] ;
wire \u_lsu.pmem[1317] ;
wire \u_lsu.pmem[1318] ;
wire \u_lsu.pmem[1319] ;
wire \u_lsu.pmem[1320] ;
wire \u_lsu.pmem[1321] ;
wire \u_lsu.pmem[1322] ;
wire \u_lsu.pmem[1323] ;
wire \u_lsu.pmem[1324] ;
wire \u_lsu.pmem[1325] ;
wire \u_lsu.pmem[1326] ;
wire \u_lsu.pmem[1327] ;
wire \u_lsu.pmem[1328] ;
wire \u_lsu.pmem[1329] ;
wire \u_lsu.pmem[1330] ;
wire \u_lsu.pmem[1331] ;
wire \u_lsu.pmem[1332] ;
wire \u_lsu.pmem[1333] ;
wire \u_lsu.pmem[1334] ;
wire \u_lsu.pmem[1335] ;
wire \u_lsu.pmem[1336] ;
wire \u_lsu.pmem[1337] ;
wire \u_lsu.pmem[1338] ;
wire \u_lsu.pmem[1339] ;
wire \u_lsu.pmem[1340] ;
wire \u_lsu.pmem[1341] ;
wire \u_lsu.pmem[1342] ;
wire \u_lsu.pmem[1343] ;
wire \u_lsu.pmem[1344] ;
wire \u_lsu.pmem[1345] ;
wire \u_lsu.pmem[1346] ;
wire \u_lsu.pmem[1347] ;
wire \u_lsu.pmem[1348] ;
wire \u_lsu.pmem[1349] ;
wire \u_lsu.pmem[1350] ;
wire \u_lsu.pmem[1351] ;
wire \u_lsu.pmem[1352] ;
wire \u_lsu.pmem[1353] ;
wire \u_lsu.pmem[1354] ;
wire \u_lsu.pmem[1355] ;
wire \u_lsu.pmem[1356] ;
wire \u_lsu.pmem[1357] ;
wire \u_lsu.pmem[1358] ;
wire \u_lsu.pmem[1359] ;
wire \u_lsu.pmem[1360] ;
wire \u_lsu.pmem[1361] ;
wire \u_lsu.pmem[1362] ;
wire \u_lsu.pmem[1363] ;
wire \u_lsu.pmem[1364] ;
wire \u_lsu.pmem[1365] ;
wire \u_lsu.pmem[1366] ;
wire \u_lsu.pmem[1367] ;
wire \u_lsu.pmem[1368] ;
wire \u_lsu.pmem[1369] ;
wire \u_lsu.pmem[1370] ;
wire \u_lsu.pmem[1371] ;
wire \u_lsu.pmem[1372] ;
wire \u_lsu.pmem[1373] ;
wire \u_lsu.pmem[1374] ;
wire \u_lsu.pmem[1375] ;
wire \u_lsu.pmem[1376] ;
wire \u_lsu.pmem[1377] ;
wire \u_lsu.pmem[1378] ;
wire \u_lsu.pmem[1379] ;
wire \u_lsu.pmem[1380] ;
wire \u_lsu.pmem[1381] ;
wire \u_lsu.pmem[1382] ;
wire \u_lsu.pmem[1383] ;
wire \u_lsu.pmem[1384] ;
wire \u_lsu.pmem[1385] ;
wire \u_lsu.pmem[1386] ;
wire \u_lsu.pmem[1387] ;
wire \u_lsu.pmem[1388] ;
wire \u_lsu.pmem[1389] ;
wire \u_lsu.pmem[1390] ;
wire \u_lsu.pmem[1391] ;
wire \u_lsu.pmem[1392] ;
wire \u_lsu.pmem[1393] ;
wire \u_lsu.pmem[1394] ;
wire \u_lsu.pmem[1395] ;
wire \u_lsu.pmem[1396] ;
wire \u_lsu.pmem[1397] ;
wire \u_lsu.pmem[1398] ;
wire \u_lsu.pmem[1399] ;
wire \u_lsu.pmem[1400] ;
wire \u_lsu.pmem[1401] ;
wire \u_lsu.pmem[1402] ;
wire \u_lsu.pmem[1403] ;
wire \u_lsu.pmem[1404] ;
wire \u_lsu.pmem[1405] ;
wire \u_lsu.pmem[1406] ;
wire \u_lsu.pmem[1407] ;
wire \u_lsu.pmem[1408] ;
wire \u_lsu.pmem[1409] ;
wire \u_lsu.pmem[1410] ;
wire \u_lsu.pmem[1411] ;
wire \u_lsu.pmem[1412] ;
wire \u_lsu.pmem[1413] ;
wire \u_lsu.pmem[1414] ;
wire \u_lsu.pmem[1415] ;
wire \u_lsu.pmem[1416] ;
wire \u_lsu.pmem[1417] ;
wire \u_lsu.pmem[1418] ;
wire \u_lsu.pmem[1419] ;
wire \u_lsu.pmem[1420] ;
wire \u_lsu.pmem[1421] ;
wire \u_lsu.pmem[1422] ;
wire \u_lsu.pmem[1423] ;
wire \u_lsu.pmem[1424] ;
wire \u_lsu.pmem[1425] ;
wire \u_lsu.pmem[1426] ;
wire \u_lsu.pmem[1427] ;
wire \u_lsu.pmem[1428] ;
wire \u_lsu.pmem[1429] ;
wire \u_lsu.pmem[1430] ;
wire \u_lsu.pmem[1431] ;
wire \u_lsu.pmem[1432] ;
wire \u_lsu.pmem[1433] ;
wire \u_lsu.pmem[1434] ;
wire \u_lsu.pmem[1435] ;
wire \u_lsu.pmem[1436] ;
wire \u_lsu.pmem[1437] ;
wire \u_lsu.pmem[1438] ;
wire \u_lsu.pmem[1439] ;
wire \u_lsu.pmem[1440] ;
wire \u_lsu.pmem[1441] ;
wire \u_lsu.pmem[1442] ;
wire \u_lsu.pmem[1443] ;
wire \u_lsu.pmem[1444] ;
wire \u_lsu.pmem[1445] ;
wire \u_lsu.pmem[1446] ;
wire \u_lsu.pmem[1447] ;
wire \u_lsu.pmem[1448] ;
wire \u_lsu.pmem[1449] ;
wire \u_lsu.pmem[1450] ;
wire \u_lsu.pmem[1451] ;
wire \u_lsu.pmem[1452] ;
wire \u_lsu.pmem[1453] ;
wire \u_lsu.pmem[1454] ;
wire \u_lsu.pmem[1455] ;
wire \u_lsu.pmem[1456] ;
wire \u_lsu.pmem[1457] ;
wire \u_lsu.pmem[1458] ;
wire \u_lsu.pmem[1459] ;
wire \u_lsu.pmem[1460] ;
wire \u_lsu.pmem[1461] ;
wire \u_lsu.pmem[1462] ;
wire \u_lsu.pmem[1463] ;
wire \u_lsu.pmem[1464] ;
wire \u_lsu.pmem[1465] ;
wire \u_lsu.pmem[1466] ;
wire \u_lsu.pmem[1467] ;
wire \u_lsu.pmem[1468] ;
wire \u_lsu.pmem[1469] ;
wire \u_lsu.pmem[1470] ;
wire \u_lsu.pmem[1471] ;
wire \u_lsu.pmem[1472] ;
wire \u_lsu.pmem[1473] ;
wire \u_lsu.pmem[1474] ;
wire \u_lsu.pmem[1475] ;
wire \u_lsu.pmem[1476] ;
wire \u_lsu.pmem[1477] ;
wire \u_lsu.pmem[1478] ;
wire \u_lsu.pmem[1479] ;
wire \u_lsu.pmem[1480] ;
wire \u_lsu.pmem[1481] ;
wire \u_lsu.pmem[1482] ;
wire \u_lsu.pmem[1483] ;
wire \u_lsu.pmem[1484] ;
wire \u_lsu.pmem[1485] ;
wire \u_lsu.pmem[1486] ;
wire \u_lsu.pmem[1487] ;
wire \u_lsu.pmem[1488] ;
wire \u_lsu.pmem[1489] ;
wire \u_lsu.pmem[1490] ;
wire \u_lsu.pmem[1491] ;
wire \u_lsu.pmem[1492] ;
wire \u_lsu.pmem[1493] ;
wire \u_lsu.pmem[1494] ;
wire \u_lsu.pmem[1495] ;
wire \u_lsu.pmem[1496] ;
wire \u_lsu.pmem[1497] ;
wire \u_lsu.pmem[1498] ;
wire \u_lsu.pmem[1499] ;
wire \u_lsu.pmem[1500] ;
wire \u_lsu.pmem[1501] ;
wire \u_lsu.pmem[1502] ;
wire \u_lsu.pmem[1503] ;
wire \u_lsu.pmem[1504] ;
wire \u_lsu.pmem[1505] ;
wire \u_lsu.pmem[1506] ;
wire \u_lsu.pmem[1507] ;
wire \u_lsu.pmem[1508] ;
wire \u_lsu.pmem[1509] ;
wire \u_lsu.pmem[1510] ;
wire \u_lsu.pmem[1511] ;
wire \u_lsu.pmem[1512] ;
wire \u_lsu.pmem[1513] ;
wire \u_lsu.pmem[1514] ;
wire \u_lsu.pmem[1515] ;
wire \u_lsu.pmem[1516] ;
wire \u_lsu.pmem[1517] ;
wire \u_lsu.pmem[1518] ;
wire \u_lsu.pmem[1519] ;
wire \u_lsu.pmem[1520] ;
wire \u_lsu.pmem[1521] ;
wire \u_lsu.pmem[1522] ;
wire \u_lsu.pmem[1523] ;
wire \u_lsu.pmem[1524] ;
wire \u_lsu.pmem[1525] ;
wire \u_lsu.pmem[1526] ;
wire \u_lsu.pmem[1527] ;
wire \u_lsu.pmem[1528] ;
wire \u_lsu.pmem[1529] ;
wire \u_lsu.pmem[1530] ;
wire \u_lsu.pmem[1531] ;
wire \u_lsu.pmem[1532] ;
wire \u_lsu.pmem[1533] ;
wire \u_lsu.pmem[1534] ;
wire \u_lsu.pmem[1535] ;
wire \u_lsu.pmem[1536] ;
wire \u_lsu.pmem[1537] ;
wire \u_lsu.pmem[1538] ;
wire \u_lsu.pmem[1539] ;
wire \u_lsu.pmem[1540] ;
wire \u_lsu.pmem[1541] ;
wire \u_lsu.pmem[1542] ;
wire \u_lsu.pmem[1543] ;
wire \u_lsu.pmem[1544] ;
wire \u_lsu.pmem[1545] ;
wire \u_lsu.pmem[1546] ;
wire \u_lsu.pmem[1547] ;
wire \u_lsu.pmem[1548] ;
wire \u_lsu.pmem[1549] ;
wire \u_lsu.pmem[1550] ;
wire \u_lsu.pmem[1551] ;
wire \u_lsu.pmem[1552] ;
wire \u_lsu.pmem[1553] ;
wire \u_lsu.pmem[1554] ;
wire \u_lsu.pmem[1555] ;
wire \u_lsu.pmem[1556] ;
wire \u_lsu.pmem[1557] ;
wire \u_lsu.pmem[1558] ;
wire \u_lsu.pmem[1559] ;
wire \u_lsu.pmem[1560] ;
wire \u_lsu.pmem[1561] ;
wire \u_lsu.pmem[1562] ;
wire \u_lsu.pmem[1563] ;
wire \u_lsu.pmem[1564] ;
wire \u_lsu.pmem[1565] ;
wire \u_lsu.pmem[1566] ;
wire \u_lsu.pmem[1567] ;
wire \u_lsu.pmem[1568] ;
wire \u_lsu.pmem[1569] ;
wire \u_lsu.pmem[1570] ;
wire \u_lsu.pmem[1571] ;
wire \u_lsu.pmem[1572] ;
wire \u_lsu.pmem[1573] ;
wire \u_lsu.pmem[1574] ;
wire \u_lsu.pmem[1575] ;
wire \u_lsu.pmem[1576] ;
wire \u_lsu.pmem[1577] ;
wire \u_lsu.pmem[1578] ;
wire \u_lsu.pmem[1579] ;
wire \u_lsu.pmem[1580] ;
wire \u_lsu.pmem[1581] ;
wire \u_lsu.pmem[1582] ;
wire \u_lsu.pmem[1583] ;
wire \u_lsu.pmem[1584] ;
wire \u_lsu.pmem[1585] ;
wire \u_lsu.pmem[1586] ;
wire \u_lsu.pmem[1587] ;
wire \u_lsu.pmem[1588] ;
wire \u_lsu.pmem[1589] ;
wire \u_lsu.pmem[1590] ;
wire \u_lsu.pmem[1591] ;
wire \u_lsu.pmem[1592] ;
wire \u_lsu.pmem[1593] ;
wire \u_lsu.pmem[1594] ;
wire \u_lsu.pmem[1595] ;
wire \u_lsu.pmem[1596] ;
wire \u_lsu.pmem[1597] ;
wire \u_lsu.pmem[1598] ;
wire \u_lsu.pmem[1599] ;
wire \u_lsu.pmem[1600] ;
wire \u_lsu.pmem[1601] ;
wire \u_lsu.pmem[1602] ;
wire \u_lsu.pmem[1603] ;
wire \u_lsu.pmem[1604] ;
wire \u_lsu.pmem[1605] ;
wire \u_lsu.pmem[1606] ;
wire \u_lsu.pmem[1607] ;
wire \u_lsu.pmem[1608] ;
wire \u_lsu.pmem[1609] ;
wire \u_lsu.pmem[1610] ;
wire \u_lsu.pmem[1611] ;
wire \u_lsu.pmem[1612] ;
wire \u_lsu.pmem[1613] ;
wire \u_lsu.pmem[1614] ;
wire \u_lsu.pmem[1615] ;
wire \u_lsu.pmem[1616] ;
wire \u_lsu.pmem[1617] ;
wire \u_lsu.pmem[1618] ;
wire \u_lsu.pmem[1619] ;
wire \u_lsu.pmem[1620] ;
wire \u_lsu.pmem[1621] ;
wire \u_lsu.pmem[1622] ;
wire \u_lsu.pmem[1623] ;
wire \u_lsu.pmem[1624] ;
wire \u_lsu.pmem[1625] ;
wire \u_lsu.pmem[1626] ;
wire \u_lsu.pmem[1627] ;
wire \u_lsu.pmem[1628] ;
wire \u_lsu.pmem[1629] ;
wire \u_lsu.pmem[1630] ;
wire \u_lsu.pmem[1631] ;
wire \u_lsu.pmem[1632] ;
wire \u_lsu.pmem[1633] ;
wire \u_lsu.pmem[1634] ;
wire \u_lsu.pmem[1635] ;
wire \u_lsu.pmem[1636] ;
wire \u_lsu.pmem[1637] ;
wire \u_lsu.pmem[1638] ;
wire \u_lsu.pmem[1639] ;
wire \u_lsu.pmem[1640] ;
wire \u_lsu.pmem[1641] ;
wire \u_lsu.pmem[1642] ;
wire \u_lsu.pmem[1643] ;
wire \u_lsu.pmem[1644] ;
wire \u_lsu.pmem[1645] ;
wire \u_lsu.pmem[1646] ;
wire \u_lsu.pmem[1647] ;
wire \u_lsu.pmem[1648] ;
wire \u_lsu.pmem[1649] ;
wire \u_lsu.pmem[1650] ;
wire \u_lsu.pmem[1651] ;
wire \u_lsu.pmem[1652] ;
wire \u_lsu.pmem[1653] ;
wire \u_lsu.pmem[1654] ;
wire \u_lsu.pmem[1655] ;
wire \u_lsu.pmem[1656] ;
wire \u_lsu.pmem[1657] ;
wire \u_lsu.pmem[1658] ;
wire \u_lsu.pmem[1659] ;
wire \u_lsu.pmem[1660] ;
wire \u_lsu.pmem[1661] ;
wire \u_lsu.pmem[1662] ;
wire \u_lsu.pmem[1663] ;
wire \u_lsu.pmem[1664] ;
wire \u_lsu.pmem[1665] ;
wire \u_lsu.pmem[1666] ;
wire \u_lsu.pmem[1667] ;
wire \u_lsu.pmem[1668] ;
wire \u_lsu.pmem[1669] ;
wire \u_lsu.pmem[1670] ;
wire \u_lsu.pmem[1671] ;
wire \u_lsu.pmem[1672] ;
wire \u_lsu.pmem[1673] ;
wire \u_lsu.pmem[1674] ;
wire \u_lsu.pmem[1675] ;
wire \u_lsu.pmem[1676] ;
wire \u_lsu.pmem[1677] ;
wire \u_lsu.pmem[1678] ;
wire \u_lsu.pmem[1679] ;
wire \u_lsu.pmem[1680] ;
wire \u_lsu.pmem[1681] ;
wire \u_lsu.pmem[1682] ;
wire \u_lsu.pmem[1683] ;
wire \u_lsu.pmem[1684] ;
wire \u_lsu.pmem[1685] ;
wire \u_lsu.pmem[1686] ;
wire \u_lsu.pmem[1687] ;
wire \u_lsu.pmem[1688] ;
wire \u_lsu.pmem[1689] ;
wire \u_lsu.pmem[1690] ;
wire \u_lsu.pmem[1691] ;
wire \u_lsu.pmem[1692] ;
wire \u_lsu.pmem[1693] ;
wire \u_lsu.pmem[1694] ;
wire \u_lsu.pmem[1695] ;
wire \u_lsu.pmem[1696] ;
wire \u_lsu.pmem[1697] ;
wire \u_lsu.pmem[1698] ;
wire \u_lsu.pmem[1699] ;
wire \u_lsu.pmem[1700] ;
wire \u_lsu.pmem[1701] ;
wire \u_lsu.pmem[1702] ;
wire \u_lsu.pmem[1703] ;
wire \u_lsu.pmem[1704] ;
wire \u_lsu.pmem[1705] ;
wire \u_lsu.pmem[1706] ;
wire \u_lsu.pmem[1707] ;
wire \u_lsu.pmem[1708] ;
wire \u_lsu.pmem[1709] ;
wire \u_lsu.pmem[1710] ;
wire \u_lsu.pmem[1711] ;
wire \u_lsu.pmem[1712] ;
wire \u_lsu.pmem[1713] ;
wire \u_lsu.pmem[1714] ;
wire \u_lsu.pmem[1715] ;
wire \u_lsu.pmem[1716] ;
wire \u_lsu.pmem[1717] ;
wire \u_lsu.pmem[1718] ;
wire \u_lsu.pmem[1719] ;
wire \u_lsu.pmem[1720] ;
wire \u_lsu.pmem[1721] ;
wire \u_lsu.pmem[1722] ;
wire \u_lsu.pmem[1723] ;
wire \u_lsu.pmem[1724] ;
wire \u_lsu.pmem[1725] ;
wire \u_lsu.pmem[1726] ;
wire \u_lsu.pmem[1727] ;
wire \u_lsu.pmem[1728] ;
wire \u_lsu.pmem[1729] ;
wire \u_lsu.pmem[1730] ;
wire \u_lsu.pmem[1731] ;
wire \u_lsu.pmem[1732] ;
wire \u_lsu.pmem[1733] ;
wire \u_lsu.pmem[1734] ;
wire \u_lsu.pmem[1735] ;
wire \u_lsu.pmem[1736] ;
wire \u_lsu.pmem[1737] ;
wire \u_lsu.pmem[1738] ;
wire \u_lsu.pmem[1739] ;
wire \u_lsu.pmem[1740] ;
wire \u_lsu.pmem[1741] ;
wire \u_lsu.pmem[1742] ;
wire \u_lsu.pmem[1743] ;
wire \u_lsu.pmem[1744] ;
wire \u_lsu.pmem[1745] ;
wire \u_lsu.pmem[1746] ;
wire \u_lsu.pmem[1747] ;
wire \u_lsu.pmem[1748] ;
wire \u_lsu.pmem[1749] ;
wire \u_lsu.pmem[1750] ;
wire \u_lsu.pmem[1751] ;
wire \u_lsu.pmem[1752] ;
wire \u_lsu.pmem[1753] ;
wire \u_lsu.pmem[1754] ;
wire \u_lsu.pmem[1755] ;
wire \u_lsu.pmem[1756] ;
wire \u_lsu.pmem[1757] ;
wire \u_lsu.pmem[1758] ;
wire \u_lsu.pmem[1759] ;
wire \u_lsu.pmem[1760] ;
wire \u_lsu.pmem[1761] ;
wire \u_lsu.pmem[1762] ;
wire \u_lsu.pmem[1763] ;
wire \u_lsu.pmem[1764] ;
wire \u_lsu.pmem[1765] ;
wire \u_lsu.pmem[1766] ;
wire \u_lsu.pmem[1767] ;
wire \u_lsu.pmem[1768] ;
wire \u_lsu.pmem[1769] ;
wire \u_lsu.pmem[1770] ;
wire \u_lsu.pmem[1771] ;
wire \u_lsu.pmem[1772] ;
wire \u_lsu.pmem[1773] ;
wire \u_lsu.pmem[1774] ;
wire \u_lsu.pmem[1775] ;
wire \u_lsu.pmem[1776] ;
wire \u_lsu.pmem[1777] ;
wire \u_lsu.pmem[1778] ;
wire \u_lsu.pmem[1779] ;
wire \u_lsu.pmem[1780] ;
wire \u_lsu.pmem[1781] ;
wire \u_lsu.pmem[1782] ;
wire \u_lsu.pmem[1783] ;
wire \u_lsu.pmem[1784] ;
wire \u_lsu.pmem[1785] ;
wire \u_lsu.pmem[1786] ;
wire \u_lsu.pmem[1787] ;
wire \u_lsu.pmem[1788] ;
wire \u_lsu.pmem[1789] ;
wire \u_lsu.pmem[1790] ;
wire \u_lsu.pmem[1791] ;
wire \u_lsu.pmem[1792] ;
wire \u_lsu.pmem[1793] ;
wire \u_lsu.pmem[1794] ;
wire \u_lsu.pmem[1795] ;
wire \u_lsu.pmem[1796] ;
wire \u_lsu.pmem[1797] ;
wire \u_lsu.pmem[1798] ;
wire \u_lsu.pmem[1799] ;
wire \u_lsu.pmem[1800] ;
wire \u_lsu.pmem[1801] ;
wire \u_lsu.pmem[1802] ;
wire \u_lsu.pmem[1803] ;
wire \u_lsu.pmem[1804] ;
wire \u_lsu.pmem[1805] ;
wire \u_lsu.pmem[1806] ;
wire \u_lsu.pmem[1807] ;
wire \u_lsu.pmem[1808] ;
wire \u_lsu.pmem[1809] ;
wire \u_lsu.pmem[1810] ;
wire \u_lsu.pmem[1811] ;
wire \u_lsu.pmem[1812] ;
wire \u_lsu.pmem[1813] ;
wire \u_lsu.pmem[1814] ;
wire \u_lsu.pmem[1815] ;
wire \u_lsu.pmem[1816] ;
wire \u_lsu.pmem[1817] ;
wire \u_lsu.pmem[1818] ;
wire \u_lsu.pmem[1819] ;
wire \u_lsu.pmem[1820] ;
wire \u_lsu.pmem[1821] ;
wire \u_lsu.pmem[1822] ;
wire \u_lsu.pmem[1823] ;
wire \u_lsu.pmem[1824] ;
wire \u_lsu.pmem[1825] ;
wire \u_lsu.pmem[1826] ;
wire \u_lsu.pmem[1827] ;
wire \u_lsu.pmem[1828] ;
wire \u_lsu.pmem[1829] ;
wire \u_lsu.pmem[1830] ;
wire \u_lsu.pmem[1831] ;
wire \u_lsu.pmem[1832] ;
wire \u_lsu.pmem[1833] ;
wire \u_lsu.pmem[1834] ;
wire \u_lsu.pmem[1835] ;
wire \u_lsu.pmem[1836] ;
wire \u_lsu.pmem[1837] ;
wire \u_lsu.pmem[1838] ;
wire \u_lsu.pmem[1839] ;
wire \u_lsu.pmem[1840] ;
wire \u_lsu.pmem[1841] ;
wire \u_lsu.pmem[1842] ;
wire \u_lsu.pmem[1843] ;
wire \u_lsu.pmem[1844] ;
wire \u_lsu.pmem[1845] ;
wire \u_lsu.pmem[1846] ;
wire \u_lsu.pmem[1847] ;
wire \u_lsu.pmem[1848] ;
wire \u_lsu.pmem[1849] ;
wire \u_lsu.pmem[1850] ;
wire \u_lsu.pmem[1851] ;
wire \u_lsu.pmem[1852] ;
wire \u_lsu.pmem[1853] ;
wire \u_lsu.pmem[1854] ;
wire \u_lsu.pmem[1855] ;
wire \u_lsu.pmem[1856] ;
wire \u_lsu.pmem[1857] ;
wire \u_lsu.pmem[1858] ;
wire \u_lsu.pmem[1859] ;
wire \u_lsu.pmem[1860] ;
wire \u_lsu.pmem[1861] ;
wire \u_lsu.pmem[1862] ;
wire \u_lsu.pmem[1863] ;
wire \u_lsu.pmem[1864] ;
wire \u_lsu.pmem[1865] ;
wire \u_lsu.pmem[1866] ;
wire \u_lsu.pmem[1867] ;
wire \u_lsu.pmem[1868] ;
wire \u_lsu.pmem[1869] ;
wire \u_lsu.pmem[1870] ;
wire \u_lsu.pmem[1871] ;
wire \u_lsu.pmem[1872] ;
wire \u_lsu.pmem[1873] ;
wire \u_lsu.pmem[1874] ;
wire \u_lsu.pmem[1875] ;
wire \u_lsu.pmem[1876] ;
wire \u_lsu.pmem[1877] ;
wire \u_lsu.pmem[1878] ;
wire \u_lsu.pmem[1879] ;
wire \u_lsu.pmem[1880] ;
wire \u_lsu.pmem[1881] ;
wire \u_lsu.pmem[1882] ;
wire \u_lsu.pmem[1883] ;
wire \u_lsu.pmem[1884] ;
wire \u_lsu.pmem[1885] ;
wire \u_lsu.pmem[1886] ;
wire \u_lsu.pmem[1887] ;
wire \u_lsu.pmem[1888] ;
wire \u_lsu.pmem[1889] ;
wire \u_lsu.pmem[1890] ;
wire \u_lsu.pmem[1891] ;
wire \u_lsu.pmem[1892] ;
wire \u_lsu.pmem[1893] ;
wire \u_lsu.pmem[1894] ;
wire \u_lsu.pmem[1895] ;
wire \u_lsu.pmem[1896] ;
wire \u_lsu.pmem[1897] ;
wire \u_lsu.pmem[1898] ;
wire \u_lsu.pmem[1899] ;
wire \u_lsu.pmem[1900] ;
wire \u_lsu.pmem[1901] ;
wire \u_lsu.pmem[1902] ;
wire \u_lsu.pmem[1903] ;
wire \u_lsu.pmem[1904] ;
wire \u_lsu.pmem[1905] ;
wire \u_lsu.pmem[1906] ;
wire \u_lsu.pmem[1907] ;
wire \u_lsu.pmem[1908] ;
wire \u_lsu.pmem[1909] ;
wire \u_lsu.pmem[1910] ;
wire \u_lsu.pmem[1911] ;
wire \u_lsu.pmem[1912] ;
wire \u_lsu.pmem[1913] ;
wire \u_lsu.pmem[1914] ;
wire \u_lsu.pmem[1915] ;
wire \u_lsu.pmem[1916] ;
wire \u_lsu.pmem[1917] ;
wire \u_lsu.pmem[1918] ;
wire \u_lsu.pmem[1919] ;
wire \u_lsu.pmem[1920] ;
wire \u_lsu.pmem[1921] ;
wire \u_lsu.pmem[1922] ;
wire \u_lsu.pmem[1923] ;
wire \u_lsu.pmem[1924] ;
wire \u_lsu.pmem[1925] ;
wire \u_lsu.pmem[1926] ;
wire \u_lsu.pmem[1927] ;
wire \u_lsu.pmem[1928] ;
wire \u_lsu.pmem[1929] ;
wire \u_lsu.pmem[1930] ;
wire \u_lsu.pmem[1931] ;
wire \u_lsu.pmem[1932] ;
wire \u_lsu.pmem[1933] ;
wire \u_lsu.pmem[1934] ;
wire \u_lsu.pmem[1935] ;
wire \u_lsu.pmem[1936] ;
wire \u_lsu.pmem[1937] ;
wire \u_lsu.pmem[1938] ;
wire \u_lsu.pmem[1939] ;
wire \u_lsu.pmem[1940] ;
wire \u_lsu.pmem[1941] ;
wire \u_lsu.pmem[1942] ;
wire \u_lsu.pmem[1943] ;
wire \u_lsu.pmem[1944] ;
wire \u_lsu.pmem[1945] ;
wire \u_lsu.pmem[1946] ;
wire \u_lsu.pmem[1947] ;
wire \u_lsu.pmem[1948] ;
wire \u_lsu.pmem[1949] ;
wire \u_lsu.pmem[1950] ;
wire \u_lsu.pmem[1951] ;
wire \u_lsu.pmem[1952] ;
wire \u_lsu.pmem[1953] ;
wire \u_lsu.pmem[1954] ;
wire \u_lsu.pmem[1955] ;
wire \u_lsu.pmem[1956] ;
wire \u_lsu.pmem[1957] ;
wire \u_lsu.pmem[1958] ;
wire \u_lsu.pmem[1959] ;
wire \u_lsu.pmem[1960] ;
wire \u_lsu.pmem[1961] ;
wire \u_lsu.pmem[1962] ;
wire \u_lsu.pmem[1963] ;
wire \u_lsu.pmem[1964] ;
wire \u_lsu.pmem[1965] ;
wire \u_lsu.pmem[1966] ;
wire \u_lsu.pmem[1967] ;
wire \u_lsu.pmem[1968] ;
wire \u_lsu.pmem[1969] ;
wire \u_lsu.pmem[1970] ;
wire \u_lsu.pmem[1971] ;
wire \u_lsu.pmem[1972] ;
wire \u_lsu.pmem[1973] ;
wire \u_lsu.pmem[1974] ;
wire \u_lsu.pmem[1975] ;
wire \u_lsu.pmem[1976] ;
wire \u_lsu.pmem[1977] ;
wire \u_lsu.pmem[1978] ;
wire \u_lsu.pmem[1979] ;
wire \u_lsu.pmem[1980] ;
wire \u_lsu.pmem[1981] ;
wire \u_lsu.pmem[1982] ;
wire \u_lsu.pmem[1983] ;
wire \u_lsu.pmem[1984] ;
wire \u_lsu.pmem[1985] ;
wire \u_lsu.pmem[1986] ;
wire \u_lsu.pmem[1987] ;
wire \u_lsu.pmem[1988] ;
wire \u_lsu.pmem[1989] ;
wire \u_lsu.pmem[1990] ;
wire \u_lsu.pmem[1991] ;
wire \u_lsu.pmem[1992] ;
wire \u_lsu.pmem[1993] ;
wire \u_lsu.pmem[1994] ;
wire \u_lsu.pmem[1995] ;
wire \u_lsu.pmem[1996] ;
wire \u_lsu.pmem[1997] ;
wire \u_lsu.pmem[1998] ;
wire \u_lsu.pmem[1999] ;
wire \u_lsu.pmem[2000] ;
wire \u_lsu.pmem[2001] ;
wire \u_lsu.pmem[2002] ;
wire \u_lsu.pmem[2003] ;
wire \u_lsu.pmem[2004] ;
wire \u_lsu.pmem[2005] ;
wire \u_lsu.pmem[2006] ;
wire \u_lsu.pmem[2007] ;
wire \u_lsu.pmem[2008] ;
wire \u_lsu.pmem[2009] ;
wire \u_lsu.pmem[2010] ;
wire \u_lsu.pmem[2011] ;
wire \u_lsu.pmem[2012] ;
wire \u_lsu.pmem[2013] ;
wire \u_lsu.pmem[2014] ;
wire \u_lsu.pmem[2015] ;
wire \u_lsu.pmem[2016] ;
wire \u_lsu.pmem[2017] ;
wire \u_lsu.pmem[2018] ;
wire \u_lsu.pmem[2019] ;
wire \u_lsu.pmem[2020] ;
wire \u_lsu.pmem[2021] ;
wire \u_lsu.pmem[2022] ;
wire \u_lsu.pmem[2023] ;
wire \u_lsu.pmem[2024] ;
wire \u_lsu.pmem[2025] ;
wire \u_lsu.pmem[2026] ;
wire \u_lsu.pmem[2027] ;
wire \u_lsu.pmem[2028] ;
wire \u_lsu.pmem[2029] ;
wire \u_lsu.pmem[2030] ;
wire \u_lsu.pmem[2031] ;
wire \u_lsu.pmem[2032] ;
wire \u_lsu.pmem[2033] ;
wire \u_lsu.pmem[2034] ;
wire \u_lsu.pmem[2035] ;
wire \u_lsu.pmem[2036] ;
wire \u_lsu.pmem[2037] ;
wire \u_lsu.pmem[2038] ;
wire \u_lsu.pmem[2039] ;
wire \u_lsu.pmem[2040] ;
wire \u_lsu.pmem[2041] ;
wire \u_lsu.pmem[2042] ;
wire \u_lsu.pmem[2043] ;
wire \u_lsu.pmem[2044] ;
wire \u_lsu.pmem[2045] ;
wire \u_lsu.pmem[2046] ;
wire \u_lsu.pmem[2047] ;
wire \u_lsu.pmem[2048] ;
wire \u_lsu.pmem[2049] ;
wire \u_lsu.pmem[2050] ;
wire \u_lsu.pmem[2051] ;
wire \u_lsu.pmem[2052] ;
wire \u_lsu.pmem[2053] ;
wire \u_lsu.pmem[2054] ;
wire \u_lsu.pmem[2055] ;
wire \u_lsu.pmem[2056] ;
wire \u_lsu.pmem[2057] ;
wire \u_lsu.pmem[2058] ;
wire \u_lsu.pmem[2059] ;
wire \u_lsu.pmem[2060] ;
wire \u_lsu.pmem[2061] ;
wire \u_lsu.pmem[2062] ;
wire \u_lsu.pmem[2063] ;
wire \u_lsu.pmem[2064] ;
wire \u_lsu.pmem[2065] ;
wire \u_lsu.pmem[2066] ;
wire \u_lsu.pmem[2067] ;
wire \u_lsu.pmem[2068] ;
wire \u_lsu.pmem[2069] ;
wire \u_lsu.pmem[2070] ;
wire \u_lsu.pmem[2071] ;
wire \u_lsu.pmem[2072] ;
wire \u_lsu.pmem[2073] ;
wire \u_lsu.pmem[2074] ;
wire \u_lsu.pmem[2075] ;
wire \u_lsu.pmem[2076] ;
wire \u_lsu.pmem[2077] ;
wire \u_lsu.pmem[2078] ;
wire \u_lsu.pmem[2079] ;
wire \u_lsu.pmem[2080] ;
wire \u_lsu.pmem[2081] ;
wire \u_lsu.pmem[2082] ;
wire \u_lsu.pmem[2083] ;
wire \u_lsu.pmem[2084] ;
wire \u_lsu.pmem[2085] ;
wire \u_lsu.pmem[2086] ;
wire \u_lsu.pmem[2087] ;
wire \u_lsu.pmem[2088] ;
wire \u_lsu.pmem[2089] ;
wire \u_lsu.pmem[2090] ;
wire \u_lsu.pmem[2091] ;
wire \u_lsu.pmem[2092] ;
wire \u_lsu.pmem[2093] ;
wire \u_lsu.pmem[2094] ;
wire \u_lsu.pmem[2095] ;
wire \u_lsu.pmem[2096] ;
wire \u_lsu.pmem[2097] ;
wire \u_lsu.pmem[2098] ;
wire \u_lsu.pmem[2099] ;
wire \u_lsu.pmem[2100] ;
wire \u_lsu.pmem[2101] ;
wire \u_lsu.pmem[2102] ;
wire \u_lsu.pmem[2103] ;
wire \u_lsu.pmem[2104] ;
wire \u_lsu.pmem[2105] ;
wire \u_lsu.pmem[2106] ;
wire \u_lsu.pmem[2107] ;
wire \u_lsu.pmem[2108] ;
wire \u_lsu.pmem[2109] ;
wire \u_lsu.pmem[2110] ;
wire \u_lsu.pmem[2111] ;
wire \u_lsu.pmem[2112] ;
wire \u_lsu.pmem[2113] ;
wire \u_lsu.pmem[2114] ;
wire \u_lsu.pmem[2115] ;
wire \u_lsu.pmem[2116] ;
wire \u_lsu.pmem[2117] ;
wire \u_lsu.pmem[2118] ;
wire \u_lsu.pmem[2119] ;
wire \u_lsu.pmem[2120] ;
wire \u_lsu.pmem[2121] ;
wire \u_lsu.pmem[2122] ;
wire \u_lsu.pmem[2123] ;
wire \u_lsu.pmem[2124] ;
wire \u_lsu.pmem[2125] ;
wire \u_lsu.pmem[2126] ;
wire \u_lsu.pmem[2127] ;
wire \u_lsu.pmem[2128] ;
wire \u_lsu.pmem[2129] ;
wire \u_lsu.pmem[2130] ;
wire \u_lsu.pmem[2131] ;
wire \u_lsu.pmem[2132] ;
wire \u_lsu.pmem[2133] ;
wire \u_lsu.pmem[2134] ;
wire \u_lsu.pmem[2135] ;
wire \u_lsu.pmem[2136] ;
wire \u_lsu.pmem[2137] ;
wire \u_lsu.pmem[2138] ;
wire \u_lsu.pmem[2139] ;
wire \u_lsu.pmem[2140] ;
wire \u_lsu.pmem[2141] ;
wire \u_lsu.pmem[2142] ;
wire \u_lsu.pmem[2143] ;
wire \u_lsu.pmem[2144] ;
wire \u_lsu.pmem[2145] ;
wire \u_lsu.pmem[2146] ;
wire \u_lsu.pmem[2147] ;
wire \u_lsu.pmem[2148] ;
wire \u_lsu.pmem[2149] ;
wire \u_lsu.pmem[2150] ;
wire \u_lsu.pmem[2151] ;
wire \u_lsu.pmem[2152] ;
wire \u_lsu.pmem[2153] ;
wire \u_lsu.pmem[2154] ;
wire \u_lsu.pmem[2155] ;
wire \u_lsu.pmem[2156] ;
wire \u_lsu.pmem[2157] ;
wire \u_lsu.pmem[2158] ;
wire \u_lsu.pmem[2159] ;
wire \u_lsu.pmem[2160] ;
wire \u_lsu.pmem[2161] ;
wire \u_lsu.pmem[2162] ;
wire \u_lsu.pmem[2163] ;
wire \u_lsu.pmem[2164] ;
wire \u_lsu.pmem[2165] ;
wire \u_lsu.pmem[2166] ;
wire \u_lsu.pmem[2167] ;
wire \u_lsu.pmem[2168] ;
wire \u_lsu.pmem[2169] ;
wire \u_lsu.pmem[2170] ;
wire \u_lsu.pmem[2171] ;
wire \u_lsu.pmem[2172] ;
wire \u_lsu.pmem[2173] ;
wire \u_lsu.pmem[2174] ;
wire \u_lsu.pmem[2175] ;
wire \u_lsu.pmem[2176] ;
wire \u_lsu.pmem[2177] ;
wire \u_lsu.pmem[2178] ;
wire \u_lsu.pmem[2179] ;
wire \u_lsu.pmem[2180] ;
wire \u_lsu.pmem[2181] ;
wire \u_lsu.pmem[2182] ;
wire \u_lsu.pmem[2183] ;
wire \u_lsu.pmem[2184] ;
wire \u_lsu.pmem[2185] ;
wire \u_lsu.pmem[2186] ;
wire \u_lsu.pmem[2187] ;
wire \u_lsu.pmem[2188] ;
wire \u_lsu.pmem[2189] ;
wire \u_lsu.pmem[2190] ;
wire \u_lsu.pmem[2191] ;
wire \u_lsu.pmem[2192] ;
wire \u_lsu.pmem[2193] ;
wire \u_lsu.pmem[2194] ;
wire \u_lsu.pmem[2195] ;
wire \u_lsu.pmem[2196] ;
wire \u_lsu.pmem[2197] ;
wire \u_lsu.pmem[2198] ;
wire \u_lsu.pmem[2199] ;
wire \u_lsu.pmem[2200] ;
wire \u_lsu.pmem[2201] ;
wire \u_lsu.pmem[2202] ;
wire \u_lsu.pmem[2203] ;
wire \u_lsu.pmem[2204] ;
wire \u_lsu.pmem[2205] ;
wire \u_lsu.pmem[2206] ;
wire \u_lsu.pmem[2207] ;
wire \u_lsu.pmem[2208] ;
wire \u_lsu.pmem[2209] ;
wire \u_lsu.pmem[2210] ;
wire \u_lsu.pmem[2211] ;
wire \u_lsu.pmem[2212] ;
wire \u_lsu.pmem[2213] ;
wire \u_lsu.pmem[2214] ;
wire \u_lsu.pmem[2215] ;
wire \u_lsu.pmem[2216] ;
wire \u_lsu.pmem[2217] ;
wire \u_lsu.pmem[2218] ;
wire \u_lsu.pmem[2219] ;
wire \u_lsu.pmem[2220] ;
wire \u_lsu.pmem[2221] ;
wire \u_lsu.pmem[2222] ;
wire \u_lsu.pmem[2223] ;
wire \u_lsu.pmem[2224] ;
wire \u_lsu.pmem[2225] ;
wire \u_lsu.pmem[2226] ;
wire \u_lsu.pmem[2227] ;
wire \u_lsu.pmem[2228] ;
wire \u_lsu.pmem[2229] ;
wire \u_lsu.pmem[2230] ;
wire \u_lsu.pmem[2231] ;
wire \u_lsu.pmem[2232] ;
wire \u_lsu.pmem[2233] ;
wire \u_lsu.pmem[2234] ;
wire \u_lsu.pmem[2235] ;
wire \u_lsu.pmem[2236] ;
wire \u_lsu.pmem[2237] ;
wire \u_lsu.pmem[2238] ;
wire \u_lsu.pmem[2239] ;
wire \u_lsu.pmem[2240] ;
wire \u_lsu.pmem[2241] ;
wire \u_lsu.pmem[2242] ;
wire \u_lsu.pmem[2243] ;
wire \u_lsu.pmem[2244] ;
wire \u_lsu.pmem[2245] ;
wire \u_lsu.pmem[2246] ;
wire \u_lsu.pmem[2247] ;
wire \u_lsu.pmem[2248] ;
wire \u_lsu.pmem[2249] ;
wire \u_lsu.pmem[2250] ;
wire \u_lsu.pmem[2251] ;
wire \u_lsu.pmem[2252] ;
wire \u_lsu.pmem[2253] ;
wire \u_lsu.pmem[2254] ;
wire \u_lsu.pmem[2255] ;
wire \u_lsu.pmem[2256] ;
wire \u_lsu.pmem[2257] ;
wire \u_lsu.pmem[2258] ;
wire \u_lsu.pmem[2259] ;
wire \u_lsu.pmem[2260] ;
wire \u_lsu.pmem[2261] ;
wire \u_lsu.pmem[2262] ;
wire \u_lsu.pmem[2263] ;
wire \u_lsu.pmem[2264] ;
wire \u_lsu.pmem[2265] ;
wire \u_lsu.pmem[2266] ;
wire \u_lsu.pmem[2267] ;
wire \u_lsu.pmem[2268] ;
wire \u_lsu.pmem[2269] ;
wire \u_lsu.pmem[2270] ;
wire \u_lsu.pmem[2271] ;
wire \u_lsu.pmem[2272] ;
wire \u_lsu.pmem[2273] ;
wire \u_lsu.pmem[2274] ;
wire \u_lsu.pmem[2275] ;
wire \u_lsu.pmem[2276] ;
wire \u_lsu.pmem[2277] ;
wire \u_lsu.pmem[2278] ;
wire \u_lsu.pmem[2279] ;
wire \u_lsu.pmem[2280] ;
wire \u_lsu.pmem[2281] ;
wire \u_lsu.pmem[2282] ;
wire \u_lsu.pmem[2283] ;
wire \u_lsu.pmem[2284] ;
wire \u_lsu.pmem[2285] ;
wire \u_lsu.pmem[2286] ;
wire \u_lsu.pmem[2287] ;
wire \u_lsu.pmem[2288] ;
wire \u_lsu.pmem[2289] ;
wire \u_lsu.pmem[2290] ;
wire \u_lsu.pmem[2291] ;
wire \u_lsu.pmem[2292] ;
wire \u_lsu.pmem[2293] ;
wire \u_lsu.pmem[2294] ;
wire \u_lsu.pmem[2295] ;
wire \u_lsu.pmem[2296] ;
wire \u_lsu.pmem[2297] ;
wire \u_lsu.pmem[2298] ;
wire \u_lsu.pmem[2299] ;
wire \u_lsu.pmem[2300] ;
wire \u_lsu.pmem[2301] ;
wire \u_lsu.pmem[2302] ;
wire \u_lsu.pmem[2303] ;
wire \u_lsu.pmem[2304] ;
wire \u_lsu.pmem[2305] ;
wire \u_lsu.pmem[2306] ;
wire \u_lsu.pmem[2307] ;
wire \u_lsu.pmem[2308] ;
wire \u_lsu.pmem[2309] ;
wire \u_lsu.pmem[2310] ;
wire \u_lsu.pmem[2311] ;
wire \u_lsu.pmem[2312] ;
wire \u_lsu.pmem[2313] ;
wire \u_lsu.pmem[2314] ;
wire \u_lsu.pmem[2315] ;
wire \u_lsu.pmem[2316] ;
wire \u_lsu.pmem[2317] ;
wire \u_lsu.pmem[2318] ;
wire \u_lsu.pmem[2319] ;
wire \u_lsu.pmem[2320] ;
wire \u_lsu.pmem[2321] ;
wire \u_lsu.pmem[2322] ;
wire \u_lsu.pmem[2323] ;
wire \u_lsu.pmem[2324] ;
wire \u_lsu.pmem[2325] ;
wire \u_lsu.pmem[2326] ;
wire \u_lsu.pmem[2327] ;
wire \u_lsu.pmem[2328] ;
wire \u_lsu.pmem[2329] ;
wire \u_lsu.pmem[2330] ;
wire \u_lsu.pmem[2331] ;
wire \u_lsu.pmem[2332] ;
wire \u_lsu.pmem[2333] ;
wire \u_lsu.pmem[2334] ;
wire \u_lsu.pmem[2335] ;
wire \u_lsu.pmem[2336] ;
wire \u_lsu.pmem[2337] ;
wire \u_lsu.pmem[2338] ;
wire \u_lsu.pmem[2339] ;
wire \u_lsu.pmem[2340] ;
wire \u_lsu.pmem[2341] ;
wire \u_lsu.pmem[2342] ;
wire \u_lsu.pmem[2343] ;
wire \u_lsu.pmem[2344] ;
wire \u_lsu.pmem[2345] ;
wire \u_lsu.pmem[2346] ;
wire \u_lsu.pmem[2347] ;
wire \u_lsu.pmem[2348] ;
wire \u_lsu.pmem[2349] ;
wire \u_lsu.pmem[2350] ;
wire \u_lsu.pmem[2351] ;
wire \u_lsu.pmem[2352] ;
wire \u_lsu.pmem[2353] ;
wire \u_lsu.pmem[2354] ;
wire \u_lsu.pmem[2355] ;
wire \u_lsu.pmem[2356] ;
wire \u_lsu.pmem[2357] ;
wire \u_lsu.pmem[2358] ;
wire \u_lsu.pmem[2359] ;
wire \u_lsu.pmem[2360] ;
wire \u_lsu.pmem[2361] ;
wire \u_lsu.pmem[2362] ;
wire \u_lsu.pmem[2363] ;
wire \u_lsu.pmem[2364] ;
wire \u_lsu.pmem[2365] ;
wire \u_lsu.pmem[2366] ;
wire \u_lsu.pmem[2367] ;
wire \u_lsu.pmem[2368] ;
wire \u_lsu.pmem[2369] ;
wire \u_lsu.pmem[2370] ;
wire \u_lsu.pmem[2371] ;
wire \u_lsu.pmem[2372] ;
wire \u_lsu.pmem[2373] ;
wire \u_lsu.pmem[2374] ;
wire \u_lsu.pmem[2375] ;
wire \u_lsu.pmem[2376] ;
wire \u_lsu.pmem[2377] ;
wire \u_lsu.pmem[2378] ;
wire \u_lsu.pmem[2379] ;
wire \u_lsu.pmem[2380] ;
wire \u_lsu.pmem[2381] ;
wire \u_lsu.pmem[2382] ;
wire \u_lsu.pmem[2383] ;
wire \u_lsu.pmem[2384] ;
wire \u_lsu.pmem[2385] ;
wire \u_lsu.pmem[2386] ;
wire \u_lsu.pmem[2387] ;
wire \u_lsu.pmem[2388] ;
wire \u_lsu.pmem[2389] ;
wire \u_lsu.pmem[2390] ;
wire \u_lsu.pmem[2391] ;
wire \u_lsu.pmem[2392] ;
wire \u_lsu.pmem[2393] ;
wire \u_lsu.pmem[2394] ;
wire \u_lsu.pmem[2395] ;
wire \u_lsu.pmem[2396] ;
wire \u_lsu.pmem[2397] ;
wire \u_lsu.pmem[2398] ;
wire \u_lsu.pmem[2399] ;
wire \u_lsu.pmem[2400] ;
wire \u_lsu.pmem[2401] ;
wire \u_lsu.pmem[2402] ;
wire \u_lsu.pmem[2403] ;
wire \u_lsu.pmem[2404] ;
wire \u_lsu.pmem[2405] ;
wire \u_lsu.pmem[2406] ;
wire \u_lsu.pmem[2407] ;
wire \u_lsu.pmem[2408] ;
wire \u_lsu.pmem[2409] ;
wire \u_lsu.pmem[2410] ;
wire \u_lsu.pmem[2411] ;
wire \u_lsu.pmem[2412] ;
wire \u_lsu.pmem[2413] ;
wire \u_lsu.pmem[2414] ;
wire \u_lsu.pmem[2415] ;
wire \u_lsu.pmem[2416] ;
wire \u_lsu.pmem[2417] ;
wire \u_lsu.pmem[2418] ;
wire \u_lsu.pmem[2419] ;
wire \u_lsu.pmem[2420] ;
wire \u_lsu.pmem[2421] ;
wire \u_lsu.pmem[2422] ;
wire \u_lsu.pmem[2423] ;
wire \u_lsu.pmem[2424] ;
wire \u_lsu.pmem[2425] ;
wire \u_lsu.pmem[2426] ;
wire \u_lsu.pmem[2427] ;
wire \u_lsu.pmem[2428] ;
wire \u_lsu.pmem[2429] ;
wire \u_lsu.pmem[2430] ;
wire \u_lsu.pmem[2431] ;
wire \u_lsu.pmem[2432] ;
wire \u_lsu.pmem[2433] ;
wire \u_lsu.pmem[2434] ;
wire \u_lsu.pmem[2435] ;
wire \u_lsu.pmem[2436] ;
wire \u_lsu.pmem[2437] ;
wire \u_lsu.pmem[2438] ;
wire \u_lsu.pmem[2439] ;
wire \u_lsu.pmem[2440] ;
wire \u_lsu.pmem[2441] ;
wire \u_lsu.pmem[2442] ;
wire \u_lsu.pmem[2443] ;
wire \u_lsu.pmem[2444] ;
wire \u_lsu.pmem[2445] ;
wire \u_lsu.pmem[2446] ;
wire \u_lsu.pmem[2447] ;
wire \u_lsu.pmem[2448] ;
wire \u_lsu.pmem[2449] ;
wire \u_lsu.pmem[2450] ;
wire \u_lsu.pmem[2451] ;
wire \u_lsu.pmem[2452] ;
wire \u_lsu.pmem[2453] ;
wire \u_lsu.pmem[2454] ;
wire \u_lsu.pmem[2455] ;
wire \u_lsu.pmem[2456] ;
wire \u_lsu.pmem[2457] ;
wire \u_lsu.pmem[2458] ;
wire \u_lsu.pmem[2459] ;
wire \u_lsu.pmem[2460] ;
wire \u_lsu.pmem[2461] ;
wire \u_lsu.pmem[2462] ;
wire \u_lsu.pmem[2463] ;
wire \u_lsu.pmem[2464] ;
wire \u_lsu.pmem[2465] ;
wire \u_lsu.pmem[2466] ;
wire \u_lsu.pmem[2467] ;
wire \u_lsu.pmem[2468] ;
wire \u_lsu.pmem[2469] ;
wire \u_lsu.pmem[2470] ;
wire \u_lsu.pmem[2471] ;
wire \u_lsu.pmem[2472] ;
wire \u_lsu.pmem[2473] ;
wire \u_lsu.pmem[2474] ;
wire \u_lsu.pmem[2475] ;
wire \u_lsu.pmem[2476] ;
wire \u_lsu.pmem[2477] ;
wire \u_lsu.pmem[2478] ;
wire \u_lsu.pmem[2479] ;
wire \u_lsu.pmem[2480] ;
wire \u_lsu.pmem[2481] ;
wire \u_lsu.pmem[2482] ;
wire \u_lsu.pmem[2483] ;
wire \u_lsu.pmem[2484] ;
wire \u_lsu.pmem[2485] ;
wire \u_lsu.pmem[2486] ;
wire \u_lsu.pmem[2487] ;
wire \u_lsu.pmem[2488] ;
wire \u_lsu.pmem[2489] ;
wire \u_lsu.pmem[2490] ;
wire \u_lsu.pmem[2491] ;
wire \u_lsu.pmem[2492] ;
wire \u_lsu.pmem[2493] ;
wire \u_lsu.pmem[2494] ;
wire \u_lsu.pmem[2495] ;
wire \u_lsu.pmem[2496] ;
wire \u_lsu.pmem[2497] ;
wire \u_lsu.pmem[2498] ;
wire \u_lsu.pmem[2499] ;
wire \u_lsu.pmem[2500] ;
wire \u_lsu.pmem[2501] ;
wire \u_lsu.pmem[2502] ;
wire \u_lsu.pmem[2503] ;
wire \u_lsu.pmem[2504] ;
wire \u_lsu.pmem[2505] ;
wire \u_lsu.pmem[2506] ;
wire \u_lsu.pmem[2507] ;
wire \u_lsu.pmem[2508] ;
wire \u_lsu.pmem[2509] ;
wire \u_lsu.pmem[2510] ;
wire \u_lsu.pmem[2511] ;
wire \u_lsu.pmem[2512] ;
wire \u_lsu.pmem[2513] ;
wire \u_lsu.pmem[2514] ;
wire \u_lsu.pmem[2515] ;
wire \u_lsu.pmem[2516] ;
wire \u_lsu.pmem[2517] ;
wire \u_lsu.pmem[2518] ;
wire \u_lsu.pmem[2519] ;
wire \u_lsu.pmem[2520] ;
wire \u_lsu.pmem[2521] ;
wire \u_lsu.pmem[2522] ;
wire \u_lsu.pmem[2523] ;
wire \u_lsu.pmem[2524] ;
wire \u_lsu.pmem[2525] ;
wire \u_lsu.pmem[2526] ;
wire \u_lsu.pmem[2527] ;
wire \u_lsu.pmem[2528] ;
wire \u_lsu.pmem[2529] ;
wire \u_lsu.pmem[2530] ;
wire \u_lsu.pmem[2531] ;
wire \u_lsu.pmem[2532] ;
wire \u_lsu.pmem[2533] ;
wire \u_lsu.pmem[2534] ;
wire \u_lsu.pmem[2535] ;
wire \u_lsu.pmem[2536] ;
wire \u_lsu.pmem[2537] ;
wire \u_lsu.pmem[2538] ;
wire \u_lsu.pmem[2539] ;
wire \u_lsu.pmem[2540] ;
wire \u_lsu.pmem[2541] ;
wire \u_lsu.pmem[2542] ;
wire \u_lsu.pmem[2543] ;
wire \u_lsu.pmem[2544] ;
wire \u_lsu.pmem[2545] ;
wire \u_lsu.pmem[2546] ;
wire \u_lsu.pmem[2547] ;
wire \u_lsu.pmem[2548] ;
wire \u_lsu.pmem[2549] ;
wire \u_lsu.pmem[2550] ;
wire \u_lsu.pmem[2551] ;
wire \u_lsu.pmem[2552] ;
wire \u_lsu.pmem[2553] ;
wire \u_lsu.pmem[2554] ;
wire \u_lsu.pmem[2555] ;
wire \u_lsu.pmem[2556] ;
wire \u_lsu.pmem[2557] ;
wire \u_lsu.pmem[2558] ;
wire \u_lsu.pmem[2559] ;
wire \u_lsu.pmem[2560] ;
wire \u_lsu.pmem[2561] ;
wire \u_lsu.pmem[2562] ;
wire \u_lsu.pmem[2563] ;
wire \u_lsu.pmem[2564] ;
wire \u_lsu.pmem[2565] ;
wire \u_lsu.pmem[2566] ;
wire \u_lsu.pmem[2567] ;
wire \u_lsu.pmem[2568] ;
wire \u_lsu.pmem[2569] ;
wire \u_lsu.pmem[2570] ;
wire \u_lsu.pmem[2571] ;
wire \u_lsu.pmem[2572] ;
wire \u_lsu.pmem[2573] ;
wire \u_lsu.pmem[2574] ;
wire \u_lsu.pmem[2575] ;
wire \u_lsu.pmem[2576] ;
wire \u_lsu.pmem[2577] ;
wire \u_lsu.pmem[2578] ;
wire \u_lsu.pmem[2579] ;
wire \u_lsu.pmem[2580] ;
wire \u_lsu.pmem[2581] ;
wire \u_lsu.pmem[2582] ;
wire \u_lsu.pmem[2583] ;
wire \u_lsu.pmem[2584] ;
wire \u_lsu.pmem[2585] ;
wire \u_lsu.pmem[2586] ;
wire \u_lsu.pmem[2587] ;
wire \u_lsu.pmem[2588] ;
wire \u_lsu.pmem[2589] ;
wire \u_lsu.pmem[2590] ;
wire \u_lsu.pmem[2591] ;
wire \u_lsu.pmem[2592] ;
wire \u_lsu.pmem[2593] ;
wire \u_lsu.pmem[2594] ;
wire \u_lsu.pmem[2595] ;
wire \u_lsu.pmem[2596] ;
wire \u_lsu.pmem[2597] ;
wire \u_lsu.pmem[2598] ;
wire \u_lsu.pmem[2599] ;
wire \u_lsu.pmem[2600] ;
wire \u_lsu.pmem[2601] ;
wire \u_lsu.pmem[2602] ;
wire \u_lsu.pmem[2603] ;
wire \u_lsu.pmem[2604] ;
wire \u_lsu.pmem[2605] ;
wire \u_lsu.pmem[2606] ;
wire \u_lsu.pmem[2607] ;
wire \u_lsu.pmem[2608] ;
wire \u_lsu.pmem[2609] ;
wire \u_lsu.pmem[2610] ;
wire \u_lsu.pmem[2611] ;
wire \u_lsu.pmem[2612] ;
wire \u_lsu.pmem[2613] ;
wire \u_lsu.pmem[2614] ;
wire \u_lsu.pmem[2615] ;
wire \u_lsu.pmem[2616] ;
wire \u_lsu.pmem[2617] ;
wire \u_lsu.pmem[2618] ;
wire \u_lsu.pmem[2619] ;
wire \u_lsu.pmem[2620] ;
wire \u_lsu.pmem[2621] ;
wire \u_lsu.pmem[2622] ;
wire \u_lsu.pmem[2623] ;
wire \u_lsu.pmem[2624] ;
wire \u_lsu.pmem[2625] ;
wire \u_lsu.pmem[2626] ;
wire \u_lsu.pmem[2627] ;
wire \u_lsu.pmem[2628] ;
wire \u_lsu.pmem[2629] ;
wire \u_lsu.pmem[2630] ;
wire \u_lsu.pmem[2631] ;
wire \u_lsu.pmem[2632] ;
wire \u_lsu.pmem[2633] ;
wire \u_lsu.pmem[2634] ;
wire \u_lsu.pmem[2635] ;
wire \u_lsu.pmem[2636] ;
wire \u_lsu.pmem[2637] ;
wire \u_lsu.pmem[2638] ;
wire \u_lsu.pmem[2639] ;
wire \u_lsu.pmem[2640] ;
wire \u_lsu.pmem[2641] ;
wire \u_lsu.pmem[2642] ;
wire \u_lsu.pmem[2643] ;
wire \u_lsu.pmem[2644] ;
wire \u_lsu.pmem[2645] ;
wire \u_lsu.pmem[2646] ;
wire \u_lsu.pmem[2647] ;
wire \u_lsu.pmem[2648] ;
wire \u_lsu.pmem[2649] ;
wire \u_lsu.pmem[2650] ;
wire \u_lsu.pmem[2651] ;
wire \u_lsu.pmem[2652] ;
wire \u_lsu.pmem[2653] ;
wire \u_lsu.pmem[2654] ;
wire \u_lsu.pmem[2655] ;
wire \u_lsu.pmem[2656] ;
wire \u_lsu.pmem[2657] ;
wire \u_lsu.pmem[2658] ;
wire \u_lsu.pmem[2659] ;
wire \u_lsu.pmem[2660] ;
wire \u_lsu.pmem[2661] ;
wire \u_lsu.pmem[2662] ;
wire \u_lsu.pmem[2663] ;
wire \u_lsu.pmem[2664] ;
wire \u_lsu.pmem[2665] ;
wire \u_lsu.pmem[2666] ;
wire \u_lsu.pmem[2667] ;
wire \u_lsu.pmem[2668] ;
wire \u_lsu.pmem[2669] ;
wire \u_lsu.pmem[2670] ;
wire \u_lsu.pmem[2671] ;
wire \u_lsu.pmem[2672] ;
wire \u_lsu.pmem[2673] ;
wire \u_lsu.pmem[2674] ;
wire \u_lsu.pmem[2675] ;
wire \u_lsu.pmem[2676] ;
wire \u_lsu.pmem[2677] ;
wire \u_lsu.pmem[2678] ;
wire \u_lsu.pmem[2679] ;
wire \u_lsu.pmem[2680] ;
wire \u_lsu.pmem[2681] ;
wire \u_lsu.pmem[2682] ;
wire \u_lsu.pmem[2683] ;
wire \u_lsu.pmem[2684] ;
wire \u_lsu.pmem[2685] ;
wire \u_lsu.pmem[2686] ;
wire \u_lsu.pmem[2687] ;
wire \u_lsu.pmem[2688] ;
wire \u_lsu.pmem[2689] ;
wire \u_lsu.pmem[2690] ;
wire \u_lsu.pmem[2691] ;
wire \u_lsu.pmem[2692] ;
wire \u_lsu.pmem[2693] ;
wire \u_lsu.pmem[2694] ;
wire \u_lsu.pmem[2695] ;
wire \u_lsu.pmem[2696] ;
wire \u_lsu.pmem[2697] ;
wire \u_lsu.pmem[2698] ;
wire \u_lsu.pmem[2699] ;
wire \u_lsu.pmem[2700] ;
wire \u_lsu.pmem[2701] ;
wire \u_lsu.pmem[2702] ;
wire \u_lsu.pmem[2703] ;
wire \u_lsu.pmem[2704] ;
wire \u_lsu.pmem[2705] ;
wire \u_lsu.pmem[2706] ;
wire \u_lsu.pmem[2707] ;
wire \u_lsu.pmem[2708] ;
wire \u_lsu.pmem[2709] ;
wire \u_lsu.pmem[2710] ;
wire \u_lsu.pmem[2711] ;
wire \u_lsu.pmem[2712] ;
wire \u_lsu.pmem[2713] ;
wire \u_lsu.pmem[2714] ;
wire \u_lsu.pmem[2715] ;
wire \u_lsu.pmem[2716] ;
wire \u_lsu.pmem[2717] ;
wire \u_lsu.pmem[2718] ;
wire \u_lsu.pmem[2719] ;
wire \u_lsu.pmem[2720] ;
wire \u_lsu.pmem[2721] ;
wire \u_lsu.pmem[2722] ;
wire \u_lsu.pmem[2723] ;
wire \u_lsu.pmem[2724] ;
wire \u_lsu.pmem[2725] ;
wire \u_lsu.pmem[2726] ;
wire \u_lsu.pmem[2727] ;
wire \u_lsu.pmem[2728] ;
wire \u_lsu.pmem[2729] ;
wire \u_lsu.pmem[2730] ;
wire \u_lsu.pmem[2731] ;
wire \u_lsu.pmem[2732] ;
wire \u_lsu.pmem[2733] ;
wire \u_lsu.pmem[2734] ;
wire \u_lsu.pmem[2735] ;
wire \u_lsu.pmem[2736] ;
wire \u_lsu.pmem[2737] ;
wire \u_lsu.pmem[2738] ;
wire \u_lsu.pmem[2739] ;
wire \u_lsu.pmem[2740] ;
wire \u_lsu.pmem[2741] ;
wire \u_lsu.pmem[2742] ;
wire \u_lsu.pmem[2743] ;
wire \u_lsu.pmem[2744] ;
wire \u_lsu.pmem[2745] ;
wire \u_lsu.pmem[2746] ;
wire \u_lsu.pmem[2747] ;
wire \u_lsu.pmem[2748] ;
wire \u_lsu.pmem[2749] ;
wire \u_lsu.pmem[2750] ;
wire \u_lsu.pmem[2751] ;
wire \u_lsu.pmem[2752] ;
wire \u_lsu.pmem[2753] ;
wire \u_lsu.pmem[2754] ;
wire \u_lsu.pmem[2755] ;
wire \u_lsu.pmem[2756] ;
wire \u_lsu.pmem[2757] ;
wire \u_lsu.pmem[2758] ;
wire \u_lsu.pmem[2759] ;
wire \u_lsu.pmem[2760] ;
wire \u_lsu.pmem[2761] ;
wire \u_lsu.pmem[2762] ;
wire \u_lsu.pmem[2763] ;
wire \u_lsu.pmem[2764] ;
wire \u_lsu.pmem[2765] ;
wire \u_lsu.pmem[2766] ;
wire \u_lsu.pmem[2767] ;
wire \u_lsu.pmem[2768] ;
wire \u_lsu.pmem[2769] ;
wire \u_lsu.pmem[2770] ;
wire \u_lsu.pmem[2771] ;
wire \u_lsu.pmem[2772] ;
wire \u_lsu.pmem[2773] ;
wire \u_lsu.pmem[2774] ;
wire \u_lsu.pmem[2775] ;
wire \u_lsu.pmem[2776] ;
wire \u_lsu.pmem[2777] ;
wire \u_lsu.pmem[2778] ;
wire \u_lsu.pmem[2779] ;
wire \u_lsu.pmem[2780] ;
wire \u_lsu.pmem[2781] ;
wire \u_lsu.pmem[2782] ;
wire \u_lsu.pmem[2783] ;
wire \u_lsu.pmem[2784] ;
wire \u_lsu.pmem[2785] ;
wire \u_lsu.pmem[2786] ;
wire \u_lsu.pmem[2787] ;
wire \u_lsu.pmem[2788] ;
wire \u_lsu.pmem[2789] ;
wire \u_lsu.pmem[2790] ;
wire \u_lsu.pmem[2791] ;
wire \u_lsu.pmem[2792] ;
wire \u_lsu.pmem[2793] ;
wire \u_lsu.pmem[2794] ;
wire \u_lsu.pmem[2795] ;
wire \u_lsu.pmem[2796] ;
wire \u_lsu.pmem[2797] ;
wire \u_lsu.pmem[2798] ;
wire \u_lsu.pmem[2799] ;
wire \u_lsu.pmem[2800] ;
wire \u_lsu.pmem[2801] ;
wire \u_lsu.pmem[2802] ;
wire \u_lsu.pmem[2803] ;
wire \u_lsu.pmem[2804] ;
wire \u_lsu.pmem[2805] ;
wire \u_lsu.pmem[2806] ;
wire \u_lsu.pmem[2807] ;
wire \u_lsu.pmem[2808] ;
wire \u_lsu.pmem[2809] ;
wire \u_lsu.pmem[2810] ;
wire \u_lsu.pmem[2811] ;
wire \u_lsu.pmem[2812] ;
wire \u_lsu.pmem[2813] ;
wire \u_lsu.pmem[2814] ;
wire \u_lsu.pmem[2815] ;
wire \u_lsu.pmem[2816] ;
wire \u_lsu.pmem[2817] ;
wire \u_lsu.pmem[2818] ;
wire \u_lsu.pmem[2819] ;
wire \u_lsu.pmem[2820] ;
wire \u_lsu.pmem[2821] ;
wire \u_lsu.pmem[2822] ;
wire \u_lsu.pmem[2823] ;
wire \u_lsu.pmem[2824] ;
wire \u_lsu.pmem[2825] ;
wire \u_lsu.pmem[2826] ;
wire \u_lsu.pmem[2827] ;
wire \u_lsu.pmem[2828] ;
wire \u_lsu.pmem[2829] ;
wire \u_lsu.pmem[2830] ;
wire \u_lsu.pmem[2831] ;
wire \u_lsu.pmem[2832] ;
wire \u_lsu.pmem[2833] ;
wire \u_lsu.pmem[2834] ;
wire \u_lsu.pmem[2835] ;
wire \u_lsu.pmem[2836] ;
wire \u_lsu.pmem[2837] ;
wire \u_lsu.pmem[2838] ;
wire \u_lsu.pmem[2839] ;
wire \u_lsu.pmem[2840] ;
wire \u_lsu.pmem[2841] ;
wire \u_lsu.pmem[2842] ;
wire \u_lsu.pmem[2843] ;
wire \u_lsu.pmem[2844] ;
wire \u_lsu.pmem[2845] ;
wire \u_lsu.pmem[2846] ;
wire \u_lsu.pmem[2847] ;
wire \u_lsu.pmem[2848] ;
wire \u_lsu.pmem[2849] ;
wire \u_lsu.pmem[2850] ;
wire \u_lsu.pmem[2851] ;
wire \u_lsu.pmem[2852] ;
wire \u_lsu.pmem[2853] ;
wire \u_lsu.pmem[2854] ;
wire \u_lsu.pmem[2855] ;
wire \u_lsu.pmem[2856] ;
wire \u_lsu.pmem[2857] ;
wire \u_lsu.pmem[2858] ;
wire \u_lsu.pmem[2859] ;
wire \u_lsu.pmem[2860] ;
wire \u_lsu.pmem[2861] ;
wire \u_lsu.pmem[2862] ;
wire \u_lsu.pmem[2863] ;
wire \u_lsu.pmem[2864] ;
wire \u_lsu.pmem[2865] ;
wire \u_lsu.pmem[2866] ;
wire \u_lsu.pmem[2867] ;
wire \u_lsu.pmem[2868] ;
wire \u_lsu.pmem[2869] ;
wire \u_lsu.pmem[2870] ;
wire \u_lsu.pmem[2871] ;
wire \u_lsu.pmem[2872] ;
wire \u_lsu.pmem[2873] ;
wire \u_lsu.pmem[2874] ;
wire \u_lsu.pmem[2875] ;
wire \u_lsu.pmem[2876] ;
wire \u_lsu.pmem[2877] ;
wire \u_lsu.pmem[2878] ;
wire \u_lsu.pmem[2879] ;
wire \u_lsu.pmem[2880] ;
wire \u_lsu.pmem[2881] ;
wire \u_lsu.pmem[2882] ;
wire \u_lsu.pmem[2883] ;
wire \u_lsu.pmem[2884] ;
wire \u_lsu.pmem[2885] ;
wire \u_lsu.pmem[2886] ;
wire \u_lsu.pmem[2887] ;
wire \u_lsu.pmem[2888] ;
wire \u_lsu.pmem[2889] ;
wire \u_lsu.pmem[2890] ;
wire \u_lsu.pmem[2891] ;
wire \u_lsu.pmem[2892] ;
wire \u_lsu.pmem[2893] ;
wire \u_lsu.pmem[2894] ;
wire \u_lsu.pmem[2895] ;
wire \u_lsu.pmem[2896] ;
wire \u_lsu.pmem[2897] ;
wire \u_lsu.pmem[2898] ;
wire \u_lsu.pmem[2899] ;
wire \u_lsu.pmem[2900] ;
wire \u_lsu.pmem[2901] ;
wire \u_lsu.pmem[2902] ;
wire \u_lsu.pmem[2903] ;
wire \u_lsu.pmem[2904] ;
wire \u_lsu.pmem[2905] ;
wire \u_lsu.pmem[2906] ;
wire \u_lsu.pmem[2907] ;
wire \u_lsu.pmem[2908] ;
wire \u_lsu.pmem[2909] ;
wire \u_lsu.pmem[2910] ;
wire \u_lsu.pmem[2911] ;
wire \u_lsu.pmem[2912] ;
wire \u_lsu.pmem[2913] ;
wire \u_lsu.pmem[2914] ;
wire \u_lsu.pmem[2915] ;
wire \u_lsu.pmem[2916] ;
wire \u_lsu.pmem[2917] ;
wire \u_lsu.pmem[2918] ;
wire \u_lsu.pmem[2919] ;
wire \u_lsu.pmem[2920] ;
wire \u_lsu.pmem[2921] ;
wire \u_lsu.pmem[2922] ;
wire \u_lsu.pmem[2923] ;
wire \u_lsu.pmem[2924] ;
wire \u_lsu.pmem[2925] ;
wire \u_lsu.pmem[2926] ;
wire \u_lsu.pmem[2927] ;
wire \u_lsu.pmem[2928] ;
wire \u_lsu.pmem[2929] ;
wire \u_lsu.pmem[2930] ;
wire \u_lsu.pmem[2931] ;
wire \u_lsu.pmem[2932] ;
wire \u_lsu.pmem[2933] ;
wire \u_lsu.pmem[2934] ;
wire \u_lsu.pmem[2935] ;
wire \u_lsu.pmem[2936] ;
wire \u_lsu.pmem[2937] ;
wire \u_lsu.pmem[2938] ;
wire \u_lsu.pmem[2939] ;
wire \u_lsu.pmem[2940] ;
wire \u_lsu.pmem[2941] ;
wire \u_lsu.pmem[2942] ;
wire \u_lsu.pmem[2943] ;
wire \u_lsu.pmem[2944] ;
wire \u_lsu.pmem[2945] ;
wire \u_lsu.pmem[2946] ;
wire \u_lsu.pmem[2947] ;
wire \u_lsu.pmem[2948] ;
wire \u_lsu.pmem[2949] ;
wire \u_lsu.pmem[2950] ;
wire \u_lsu.pmem[2951] ;
wire \u_lsu.pmem[2952] ;
wire \u_lsu.pmem[2953] ;
wire \u_lsu.pmem[2954] ;
wire \u_lsu.pmem[2955] ;
wire \u_lsu.pmem[2956] ;
wire \u_lsu.pmem[2957] ;
wire \u_lsu.pmem[2958] ;
wire \u_lsu.pmem[2959] ;
wire \u_lsu.pmem[2960] ;
wire \u_lsu.pmem[2961] ;
wire \u_lsu.pmem[2962] ;
wire \u_lsu.pmem[2963] ;
wire \u_lsu.pmem[2964] ;
wire \u_lsu.pmem[2965] ;
wire \u_lsu.pmem[2966] ;
wire \u_lsu.pmem[2967] ;
wire \u_lsu.pmem[2968] ;
wire \u_lsu.pmem[2969] ;
wire \u_lsu.pmem[2970] ;
wire \u_lsu.pmem[2971] ;
wire \u_lsu.pmem[2972] ;
wire \u_lsu.pmem[2973] ;
wire \u_lsu.pmem[2974] ;
wire \u_lsu.pmem[2975] ;
wire \u_lsu.pmem[2976] ;
wire \u_lsu.pmem[2977] ;
wire \u_lsu.pmem[2978] ;
wire \u_lsu.pmem[2979] ;
wire \u_lsu.pmem[2980] ;
wire \u_lsu.pmem[2981] ;
wire \u_lsu.pmem[2982] ;
wire \u_lsu.pmem[2983] ;
wire \u_lsu.pmem[2984] ;
wire \u_lsu.pmem[2985] ;
wire \u_lsu.pmem[2986] ;
wire \u_lsu.pmem[2987] ;
wire \u_lsu.pmem[2988] ;
wire \u_lsu.pmem[2989] ;
wire \u_lsu.pmem[2990] ;
wire \u_lsu.pmem[2991] ;
wire \u_lsu.pmem[2992] ;
wire \u_lsu.pmem[2993] ;
wire \u_lsu.pmem[2994] ;
wire \u_lsu.pmem[2995] ;
wire \u_lsu.pmem[2996] ;
wire \u_lsu.pmem[2997] ;
wire \u_lsu.pmem[2998] ;
wire \u_lsu.pmem[2999] ;
wire \u_lsu.pmem[3000] ;
wire \u_lsu.pmem[3001] ;
wire \u_lsu.pmem[3002] ;
wire \u_lsu.pmem[3003] ;
wire \u_lsu.pmem[3004] ;
wire \u_lsu.pmem[3005] ;
wire \u_lsu.pmem[3006] ;
wire \u_lsu.pmem[3007] ;
wire \u_lsu.pmem[3008] ;
wire \u_lsu.pmem[3009] ;
wire \u_lsu.pmem[3010] ;
wire \u_lsu.pmem[3011] ;
wire \u_lsu.pmem[3012] ;
wire \u_lsu.pmem[3013] ;
wire \u_lsu.pmem[3014] ;
wire \u_lsu.pmem[3015] ;
wire \u_lsu.pmem[3016] ;
wire \u_lsu.pmem[3017] ;
wire \u_lsu.pmem[3018] ;
wire \u_lsu.pmem[3019] ;
wire \u_lsu.pmem[3020] ;
wire \u_lsu.pmem[3021] ;
wire \u_lsu.pmem[3022] ;
wire \u_lsu.pmem[3023] ;
wire \u_lsu.pmem[3024] ;
wire \u_lsu.pmem[3025] ;
wire \u_lsu.pmem[3026] ;
wire \u_lsu.pmem[3027] ;
wire \u_lsu.pmem[3028] ;
wire \u_lsu.pmem[3029] ;
wire \u_lsu.pmem[3030] ;
wire \u_lsu.pmem[3031] ;
wire \u_lsu.pmem[3032] ;
wire \u_lsu.pmem[3033] ;
wire \u_lsu.pmem[3034] ;
wire \u_lsu.pmem[3035] ;
wire \u_lsu.pmem[3036] ;
wire \u_lsu.pmem[3037] ;
wire \u_lsu.pmem[3038] ;
wire \u_lsu.pmem[3039] ;
wire \u_lsu.pmem[3040] ;
wire \u_lsu.pmem[3041] ;
wire \u_lsu.pmem[3042] ;
wire \u_lsu.pmem[3043] ;
wire \u_lsu.pmem[3044] ;
wire \u_lsu.pmem[3045] ;
wire \u_lsu.pmem[3046] ;
wire \u_lsu.pmem[3047] ;
wire \u_lsu.pmem[3048] ;
wire \u_lsu.pmem[3049] ;
wire \u_lsu.pmem[3050] ;
wire \u_lsu.pmem[3051] ;
wire \u_lsu.pmem[3052] ;
wire \u_lsu.pmem[3053] ;
wire \u_lsu.pmem[3054] ;
wire \u_lsu.pmem[3055] ;
wire \u_lsu.pmem[3056] ;
wire \u_lsu.pmem[3057] ;
wire \u_lsu.pmem[3058] ;
wire \u_lsu.pmem[3059] ;
wire \u_lsu.pmem[3060] ;
wire \u_lsu.pmem[3061] ;
wire \u_lsu.pmem[3062] ;
wire \u_lsu.pmem[3063] ;
wire \u_lsu.pmem[3064] ;
wire \u_lsu.pmem[3065] ;
wire \u_lsu.pmem[3066] ;
wire \u_lsu.pmem[3067] ;
wire \u_lsu.pmem[3068] ;
wire \u_lsu.pmem[3069] ;
wire \u_lsu.pmem[3070] ;
wire \u_lsu.pmem[3071] ;
wire \u_lsu.pmem[3072] ;
wire \u_lsu.pmem[3073] ;
wire \u_lsu.pmem[3074] ;
wire \u_lsu.pmem[3075] ;
wire \u_lsu.pmem[3076] ;
wire \u_lsu.pmem[3077] ;
wire \u_lsu.pmem[3078] ;
wire \u_lsu.pmem[3079] ;
wire \u_lsu.pmem[3080] ;
wire \u_lsu.pmem[3081] ;
wire \u_lsu.pmem[3082] ;
wire \u_lsu.pmem[3083] ;
wire \u_lsu.pmem[3084] ;
wire \u_lsu.pmem[3085] ;
wire \u_lsu.pmem[3086] ;
wire \u_lsu.pmem[3087] ;
wire \u_lsu.pmem[3088] ;
wire \u_lsu.pmem[3089] ;
wire \u_lsu.pmem[3090] ;
wire \u_lsu.pmem[3091] ;
wire \u_lsu.pmem[3092] ;
wire \u_lsu.pmem[3093] ;
wire \u_lsu.pmem[3094] ;
wire \u_lsu.pmem[3095] ;
wire \u_lsu.pmem[3096] ;
wire \u_lsu.pmem[3097] ;
wire \u_lsu.pmem[3098] ;
wire \u_lsu.pmem[3099] ;
wire \u_lsu.pmem[3100] ;
wire \u_lsu.pmem[3101] ;
wire \u_lsu.pmem[3102] ;
wire \u_lsu.pmem[3103] ;
wire \u_lsu.pmem[3104] ;
wire \u_lsu.pmem[3105] ;
wire \u_lsu.pmem[3106] ;
wire \u_lsu.pmem[3107] ;
wire \u_lsu.pmem[3108] ;
wire \u_lsu.pmem[3109] ;
wire \u_lsu.pmem[3110] ;
wire \u_lsu.pmem[3111] ;
wire \u_lsu.pmem[3112] ;
wire \u_lsu.pmem[3113] ;
wire \u_lsu.pmem[3114] ;
wire \u_lsu.pmem[3115] ;
wire \u_lsu.pmem[3116] ;
wire \u_lsu.pmem[3117] ;
wire \u_lsu.pmem[3118] ;
wire \u_lsu.pmem[3119] ;
wire \u_lsu.pmem[3120] ;
wire \u_lsu.pmem[3121] ;
wire \u_lsu.pmem[3122] ;
wire \u_lsu.pmem[3123] ;
wire \u_lsu.pmem[3124] ;
wire \u_lsu.pmem[3125] ;
wire \u_lsu.pmem[3126] ;
wire \u_lsu.pmem[3127] ;
wire \u_lsu.pmem[3128] ;
wire \u_lsu.pmem[3129] ;
wire \u_lsu.pmem[3130] ;
wire \u_lsu.pmem[3131] ;
wire \u_lsu.pmem[3132] ;
wire \u_lsu.pmem[3133] ;
wire \u_lsu.pmem[3134] ;
wire \u_lsu.pmem[3135] ;
wire \u_lsu.pmem[3136] ;
wire \u_lsu.pmem[3137] ;
wire \u_lsu.pmem[3138] ;
wire \u_lsu.pmem[3139] ;
wire \u_lsu.pmem[3140] ;
wire \u_lsu.pmem[3141] ;
wire \u_lsu.pmem[3142] ;
wire \u_lsu.pmem[3143] ;
wire \u_lsu.pmem[3144] ;
wire \u_lsu.pmem[3145] ;
wire \u_lsu.pmem[3146] ;
wire \u_lsu.pmem[3147] ;
wire \u_lsu.pmem[3148] ;
wire \u_lsu.pmem[3149] ;
wire \u_lsu.pmem[3150] ;
wire \u_lsu.pmem[3151] ;
wire \u_lsu.pmem[3152] ;
wire \u_lsu.pmem[3153] ;
wire \u_lsu.pmem[3154] ;
wire \u_lsu.pmem[3155] ;
wire \u_lsu.pmem[3156] ;
wire \u_lsu.pmem[3157] ;
wire \u_lsu.pmem[3158] ;
wire \u_lsu.pmem[3159] ;
wire \u_lsu.pmem[3160] ;
wire \u_lsu.pmem[3161] ;
wire \u_lsu.pmem[3162] ;
wire \u_lsu.pmem[3163] ;
wire \u_lsu.pmem[3164] ;
wire \u_lsu.pmem[3165] ;
wire \u_lsu.pmem[3166] ;
wire \u_lsu.pmem[3167] ;
wire \u_lsu.pmem[3168] ;
wire \u_lsu.pmem[3169] ;
wire \u_lsu.pmem[3170] ;
wire \u_lsu.pmem[3171] ;
wire \u_lsu.pmem[3172] ;
wire \u_lsu.pmem[3173] ;
wire \u_lsu.pmem[3174] ;
wire \u_lsu.pmem[3175] ;
wire \u_lsu.pmem[3176] ;
wire \u_lsu.pmem[3177] ;
wire \u_lsu.pmem[3178] ;
wire \u_lsu.pmem[3179] ;
wire \u_lsu.pmem[3180] ;
wire \u_lsu.pmem[3181] ;
wire \u_lsu.pmem[3182] ;
wire \u_lsu.pmem[3183] ;
wire \u_lsu.pmem[3184] ;
wire \u_lsu.pmem[3185] ;
wire \u_lsu.pmem[3186] ;
wire \u_lsu.pmem[3187] ;
wire \u_lsu.pmem[3188] ;
wire \u_lsu.pmem[3189] ;
wire \u_lsu.pmem[3190] ;
wire \u_lsu.pmem[3191] ;
wire \u_lsu.pmem[3192] ;
wire \u_lsu.pmem[3193] ;
wire \u_lsu.pmem[3194] ;
wire \u_lsu.pmem[3195] ;
wire \u_lsu.pmem[3196] ;
wire \u_lsu.pmem[3197] ;
wire \u_lsu.pmem[3198] ;
wire \u_lsu.pmem[3199] ;
wire \u_lsu.pmem[3200] ;
wire \u_lsu.pmem[3201] ;
wire \u_lsu.pmem[3202] ;
wire \u_lsu.pmem[3203] ;
wire \u_lsu.pmem[3204] ;
wire \u_lsu.pmem[3205] ;
wire \u_lsu.pmem[3206] ;
wire \u_lsu.pmem[3207] ;
wire \u_lsu.pmem[3208] ;
wire \u_lsu.pmem[3209] ;
wire \u_lsu.pmem[3210] ;
wire \u_lsu.pmem[3211] ;
wire \u_lsu.pmem[3212] ;
wire \u_lsu.pmem[3213] ;
wire \u_lsu.pmem[3214] ;
wire \u_lsu.pmem[3215] ;
wire \u_lsu.pmem[3216] ;
wire \u_lsu.pmem[3217] ;
wire \u_lsu.pmem[3218] ;
wire \u_lsu.pmem[3219] ;
wire \u_lsu.pmem[3220] ;
wire \u_lsu.pmem[3221] ;
wire \u_lsu.pmem[3222] ;
wire \u_lsu.pmem[3223] ;
wire \u_lsu.pmem[3224] ;
wire \u_lsu.pmem[3225] ;
wire \u_lsu.pmem[3226] ;
wire \u_lsu.pmem[3227] ;
wire \u_lsu.pmem[3228] ;
wire \u_lsu.pmem[3229] ;
wire \u_lsu.pmem[3230] ;
wire \u_lsu.pmem[3231] ;
wire \u_lsu.pmem[3232] ;
wire \u_lsu.pmem[3233] ;
wire \u_lsu.pmem[3234] ;
wire \u_lsu.pmem[3235] ;
wire \u_lsu.pmem[3236] ;
wire \u_lsu.pmem[3237] ;
wire \u_lsu.pmem[3238] ;
wire \u_lsu.pmem[3239] ;
wire \u_lsu.pmem[3240] ;
wire \u_lsu.pmem[3241] ;
wire \u_lsu.pmem[3242] ;
wire \u_lsu.pmem[3243] ;
wire \u_lsu.pmem[3244] ;
wire \u_lsu.pmem[3245] ;
wire \u_lsu.pmem[3246] ;
wire \u_lsu.pmem[3247] ;
wire \u_lsu.pmem[3248] ;
wire \u_lsu.pmem[3249] ;
wire \u_lsu.pmem[3250] ;
wire \u_lsu.pmem[3251] ;
wire \u_lsu.pmem[3252] ;
wire \u_lsu.pmem[3253] ;
wire \u_lsu.pmem[3254] ;
wire \u_lsu.pmem[3255] ;
wire \u_lsu.pmem[3256] ;
wire \u_lsu.pmem[3257] ;
wire \u_lsu.pmem[3258] ;
wire \u_lsu.pmem[3259] ;
wire \u_lsu.pmem[3260] ;
wire \u_lsu.pmem[3261] ;
wire \u_lsu.pmem[3262] ;
wire \u_lsu.pmem[3263] ;
wire \u_lsu.pmem[3264] ;
wire \u_lsu.pmem[3265] ;
wire \u_lsu.pmem[3266] ;
wire \u_lsu.pmem[3267] ;
wire \u_lsu.pmem[3268] ;
wire \u_lsu.pmem[3269] ;
wire \u_lsu.pmem[3270] ;
wire \u_lsu.pmem[3271] ;
wire \u_lsu.pmem[3272] ;
wire \u_lsu.pmem[3273] ;
wire \u_lsu.pmem[3274] ;
wire \u_lsu.pmem[3275] ;
wire \u_lsu.pmem[3276] ;
wire \u_lsu.pmem[3277] ;
wire \u_lsu.pmem[3278] ;
wire \u_lsu.pmem[3279] ;
wire \u_lsu.pmem[3280] ;
wire \u_lsu.pmem[3281] ;
wire \u_lsu.pmem[3282] ;
wire \u_lsu.pmem[3283] ;
wire \u_lsu.pmem[3284] ;
wire \u_lsu.pmem[3285] ;
wire \u_lsu.pmem[3286] ;
wire \u_lsu.pmem[3287] ;
wire \u_lsu.pmem[3288] ;
wire \u_lsu.pmem[3289] ;
wire \u_lsu.pmem[3290] ;
wire \u_lsu.pmem[3291] ;
wire \u_lsu.pmem[3292] ;
wire \u_lsu.pmem[3293] ;
wire \u_lsu.pmem[3294] ;
wire \u_lsu.pmem[3295] ;
wire \u_lsu.pmem[3296] ;
wire \u_lsu.pmem[3297] ;
wire \u_lsu.pmem[3298] ;
wire \u_lsu.pmem[3299] ;
wire \u_lsu.pmem[3300] ;
wire \u_lsu.pmem[3301] ;
wire \u_lsu.pmem[3302] ;
wire \u_lsu.pmem[3303] ;
wire \u_lsu.pmem[3304] ;
wire \u_lsu.pmem[3305] ;
wire \u_lsu.pmem[3306] ;
wire \u_lsu.pmem[3307] ;
wire \u_lsu.pmem[3308] ;
wire \u_lsu.pmem[3309] ;
wire \u_lsu.pmem[3310] ;
wire \u_lsu.pmem[3311] ;
wire \u_lsu.pmem[3312] ;
wire \u_lsu.pmem[3313] ;
wire \u_lsu.pmem[3314] ;
wire \u_lsu.pmem[3315] ;
wire \u_lsu.pmem[3316] ;
wire \u_lsu.pmem[3317] ;
wire \u_lsu.pmem[3318] ;
wire \u_lsu.pmem[3319] ;
wire \u_lsu.pmem[3320] ;
wire \u_lsu.pmem[3321] ;
wire \u_lsu.pmem[3322] ;
wire \u_lsu.pmem[3323] ;
wire \u_lsu.pmem[3324] ;
wire \u_lsu.pmem[3325] ;
wire \u_lsu.pmem[3326] ;
wire \u_lsu.pmem[3327] ;
wire \u_lsu.pmem[3328] ;
wire \u_lsu.pmem[3329] ;
wire \u_lsu.pmem[3330] ;
wire \u_lsu.pmem[3331] ;
wire \u_lsu.pmem[3332] ;
wire \u_lsu.pmem[3333] ;
wire \u_lsu.pmem[3334] ;
wire \u_lsu.pmem[3335] ;
wire \u_lsu.pmem[3336] ;
wire \u_lsu.pmem[3337] ;
wire \u_lsu.pmem[3338] ;
wire \u_lsu.pmem[3339] ;
wire \u_lsu.pmem[3340] ;
wire \u_lsu.pmem[3341] ;
wire \u_lsu.pmem[3342] ;
wire \u_lsu.pmem[3343] ;
wire \u_lsu.pmem[3344] ;
wire \u_lsu.pmem[3345] ;
wire \u_lsu.pmem[3346] ;
wire \u_lsu.pmem[3347] ;
wire \u_lsu.pmem[3348] ;
wire \u_lsu.pmem[3349] ;
wire \u_lsu.pmem[3350] ;
wire \u_lsu.pmem[3351] ;
wire \u_lsu.pmem[3352] ;
wire \u_lsu.pmem[3353] ;
wire \u_lsu.pmem[3354] ;
wire \u_lsu.pmem[3355] ;
wire \u_lsu.pmem[3356] ;
wire \u_lsu.pmem[3357] ;
wire \u_lsu.pmem[3358] ;
wire \u_lsu.pmem[3359] ;
wire \u_lsu.pmem[3360] ;
wire \u_lsu.pmem[3361] ;
wire \u_lsu.pmem[3362] ;
wire \u_lsu.pmem[3363] ;
wire \u_lsu.pmem[3364] ;
wire \u_lsu.pmem[3365] ;
wire \u_lsu.pmem[3366] ;
wire \u_lsu.pmem[3367] ;
wire \u_lsu.pmem[3368] ;
wire \u_lsu.pmem[3369] ;
wire \u_lsu.pmem[3370] ;
wire \u_lsu.pmem[3371] ;
wire \u_lsu.pmem[3372] ;
wire \u_lsu.pmem[3373] ;
wire \u_lsu.pmem[3374] ;
wire \u_lsu.pmem[3375] ;
wire \u_lsu.pmem[3376] ;
wire \u_lsu.pmem[3377] ;
wire \u_lsu.pmem[3378] ;
wire \u_lsu.pmem[3379] ;
wire \u_lsu.pmem[3380] ;
wire \u_lsu.pmem[3381] ;
wire \u_lsu.pmem[3382] ;
wire \u_lsu.pmem[3383] ;
wire \u_lsu.pmem[3384] ;
wire \u_lsu.pmem[3385] ;
wire \u_lsu.pmem[3386] ;
wire \u_lsu.pmem[3387] ;
wire \u_lsu.pmem[3388] ;
wire \u_lsu.pmem[3389] ;
wire \u_lsu.pmem[3390] ;
wire \u_lsu.pmem[3391] ;
wire \u_lsu.pmem[3392] ;
wire \u_lsu.pmem[3393] ;
wire \u_lsu.pmem[3394] ;
wire \u_lsu.pmem[3395] ;
wire \u_lsu.pmem[3396] ;
wire \u_lsu.pmem[3397] ;
wire \u_lsu.pmem[3398] ;
wire \u_lsu.pmem[3399] ;
wire \u_lsu.pmem[3400] ;
wire \u_lsu.pmem[3401] ;
wire \u_lsu.pmem[3402] ;
wire \u_lsu.pmem[3403] ;
wire \u_lsu.pmem[3404] ;
wire \u_lsu.pmem[3405] ;
wire \u_lsu.pmem[3406] ;
wire \u_lsu.pmem[3407] ;
wire \u_lsu.pmem[3408] ;
wire \u_lsu.pmem[3409] ;
wire \u_lsu.pmem[3410] ;
wire \u_lsu.pmem[3411] ;
wire \u_lsu.pmem[3412] ;
wire \u_lsu.pmem[3413] ;
wire \u_lsu.pmem[3414] ;
wire \u_lsu.pmem[3415] ;
wire \u_lsu.pmem[3416] ;
wire \u_lsu.pmem[3417] ;
wire \u_lsu.pmem[3418] ;
wire \u_lsu.pmem[3419] ;
wire \u_lsu.pmem[3420] ;
wire \u_lsu.pmem[3421] ;
wire \u_lsu.pmem[3422] ;
wire \u_lsu.pmem[3423] ;
wire \u_lsu.pmem[3424] ;
wire \u_lsu.pmem[3425] ;
wire \u_lsu.pmem[3426] ;
wire \u_lsu.pmem[3427] ;
wire \u_lsu.pmem[3428] ;
wire \u_lsu.pmem[3429] ;
wire \u_lsu.pmem[3430] ;
wire \u_lsu.pmem[3431] ;
wire \u_lsu.pmem[3432] ;
wire \u_lsu.pmem[3433] ;
wire \u_lsu.pmem[3434] ;
wire \u_lsu.pmem[3435] ;
wire \u_lsu.pmem[3436] ;
wire \u_lsu.pmem[3437] ;
wire \u_lsu.pmem[3438] ;
wire \u_lsu.pmem[3439] ;
wire \u_lsu.pmem[3440] ;
wire \u_lsu.pmem[3441] ;
wire \u_lsu.pmem[3442] ;
wire \u_lsu.pmem[3443] ;
wire \u_lsu.pmem[3444] ;
wire \u_lsu.pmem[3445] ;
wire \u_lsu.pmem[3446] ;
wire \u_lsu.pmem[3447] ;
wire \u_lsu.pmem[3448] ;
wire \u_lsu.pmem[3449] ;
wire \u_lsu.pmem[3450] ;
wire \u_lsu.pmem[3451] ;
wire \u_lsu.pmem[3452] ;
wire \u_lsu.pmem[3453] ;
wire \u_lsu.pmem[3454] ;
wire \u_lsu.pmem[3455] ;
wire \u_lsu.pmem[3456] ;
wire \u_lsu.pmem[3457] ;
wire \u_lsu.pmem[3458] ;
wire \u_lsu.pmem[3459] ;
wire \u_lsu.pmem[3460] ;
wire \u_lsu.pmem[3461] ;
wire \u_lsu.pmem[3462] ;
wire \u_lsu.pmem[3463] ;
wire \u_lsu.pmem[3464] ;
wire \u_lsu.pmem[3465] ;
wire \u_lsu.pmem[3466] ;
wire \u_lsu.pmem[3467] ;
wire \u_lsu.pmem[3468] ;
wire \u_lsu.pmem[3469] ;
wire \u_lsu.pmem[3470] ;
wire \u_lsu.pmem[3471] ;
wire \u_lsu.pmem[3472] ;
wire \u_lsu.pmem[3473] ;
wire \u_lsu.pmem[3474] ;
wire \u_lsu.pmem[3475] ;
wire \u_lsu.pmem[3476] ;
wire \u_lsu.pmem[3477] ;
wire \u_lsu.pmem[3478] ;
wire \u_lsu.pmem[3479] ;
wire \u_lsu.pmem[3480] ;
wire \u_lsu.pmem[3481] ;
wire \u_lsu.pmem[3482] ;
wire \u_lsu.pmem[3483] ;
wire \u_lsu.pmem[3484] ;
wire \u_lsu.pmem[3485] ;
wire \u_lsu.pmem[3486] ;
wire \u_lsu.pmem[3487] ;
wire \u_lsu.pmem[3488] ;
wire \u_lsu.pmem[3489] ;
wire \u_lsu.pmem[3490] ;
wire \u_lsu.pmem[3491] ;
wire \u_lsu.pmem[3492] ;
wire \u_lsu.pmem[3493] ;
wire \u_lsu.pmem[3494] ;
wire \u_lsu.pmem[3495] ;
wire \u_lsu.pmem[3496] ;
wire \u_lsu.pmem[3497] ;
wire \u_lsu.pmem[3498] ;
wire \u_lsu.pmem[3499] ;
wire \u_lsu.pmem[3500] ;
wire \u_lsu.pmem[3501] ;
wire \u_lsu.pmem[3502] ;
wire \u_lsu.pmem[3503] ;
wire \u_lsu.pmem[3504] ;
wire \u_lsu.pmem[3505] ;
wire \u_lsu.pmem[3506] ;
wire \u_lsu.pmem[3507] ;
wire \u_lsu.pmem[3508] ;
wire \u_lsu.pmem[3509] ;
wire \u_lsu.pmem[3510] ;
wire \u_lsu.pmem[3511] ;
wire \u_lsu.pmem[3512] ;
wire \u_lsu.pmem[3513] ;
wire \u_lsu.pmem[3514] ;
wire \u_lsu.pmem[3515] ;
wire \u_lsu.pmem[3516] ;
wire \u_lsu.pmem[3517] ;
wire \u_lsu.pmem[3518] ;
wire \u_lsu.pmem[3519] ;
wire \u_lsu.pmem[3520] ;
wire \u_lsu.pmem[3521] ;
wire \u_lsu.pmem[3522] ;
wire \u_lsu.pmem[3523] ;
wire \u_lsu.pmem[3524] ;
wire \u_lsu.pmem[3525] ;
wire \u_lsu.pmem[3526] ;
wire \u_lsu.pmem[3527] ;
wire \u_lsu.pmem[3528] ;
wire \u_lsu.pmem[3529] ;
wire \u_lsu.pmem[3530] ;
wire \u_lsu.pmem[3531] ;
wire \u_lsu.pmem[3532] ;
wire \u_lsu.pmem[3533] ;
wire \u_lsu.pmem[3534] ;
wire \u_lsu.pmem[3535] ;
wire \u_lsu.pmem[3536] ;
wire \u_lsu.pmem[3537] ;
wire \u_lsu.pmem[3538] ;
wire \u_lsu.pmem[3539] ;
wire \u_lsu.pmem[3540] ;
wire \u_lsu.pmem[3541] ;
wire \u_lsu.pmem[3542] ;
wire \u_lsu.pmem[3543] ;
wire \u_lsu.pmem[3544] ;
wire \u_lsu.pmem[3545] ;
wire \u_lsu.pmem[3546] ;
wire \u_lsu.pmem[3547] ;
wire \u_lsu.pmem[3548] ;
wire \u_lsu.pmem[3549] ;
wire \u_lsu.pmem[3550] ;
wire \u_lsu.pmem[3551] ;
wire \u_lsu.pmem[3552] ;
wire \u_lsu.pmem[3553] ;
wire \u_lsu.pmem[3554] ;
wire \u_lsu.pmem[3555] ;
wire \u_lsu.pmem[3556] ;
wire \u_lsu.pmem[3557] ;
wire \u_lsu.pmem[3558] ;
wire \u_lsu.pmem[3559] ;
wire \u_lsu.pmem[3560] ;
wire \u_lsu.pmem[3561] ;
wire \u_lsu.pmem[3562] ;
wire \u_lsu.pmem[3563] ;
wire \u_lsu.pmem[3564] ;
wire \u_lsu.pmem[3565] ;
wire \u_lsu.pmem[3566] ;
wire \u_lsu.pmem[3567] ;
wire \u_lsu.pmem[3568] ;
wire \u_lsu.pmem[3569] ;
wire \u_lsu.pmem[3570] ;
wire \u_lsu.pmem[3571] ;
wire \u_lsu.pmem[3572] ;
wire \u_lsu.pmem[3573] ;
wire \u_lsu.pmem[3574] ;
wire \u_lsu.pmem[3575] ;
wire \u_lsu.pmem[3576] ;
wire \u_lsu.pmem[3577] ;
wire \u_lsu.pmem[3578] ;
wire \u_lsu.pmem[3579] ;
wire \u_lsu.pmem[3580] ;
wire \u_lsu.pmem[3581] ;
wire \u_lsu.pmem[3582] ;
wire \u_lsu.pmem[3583] ;
wire \u_lsu.pmem[3584] ;
wire \u_lsu.pmem[3585] ;
wire \u_lsu.pmem[3586] ;
wire \u_lsu.pmem[3587] ;
wire \u_lsu.pmem[3588] ;
wire \u_lsu.pmem[3589] ;
wire \u_lsu.pmem[3590] ;
wire \u_lsu.pmem[3591] ;
wire \u_lsu.pmem[3592] ;
wire \u_lsu.pmem[3593] ;
wire \u_lsu.pmem[3594] ;
wire \u_lsu.pmem[3595] ;
wire \u_lsu.pmem[3596] ;
wire \u_lsu.pmem[3597] ;
wire \u_lsu.pmem[3598] ;
wire \u_lsu.pmem[3599] ;
wire \u_lsu.pmem[3600] ;
wire \u_lsu.pmem[3601] ;
wire \u_lsu.pmem[3602] ;
wire \u_lsu.pmem[3603] ;
wire \u_lsu.pmem[3604] ;
wire \u_lsu.pmem[3605] ;
wire \u_lsu.pmem[3606] ;
wire \u_lsu.pmem[3607] ;
wire \u_lsu.pmem[3608] ;
wire \u_lsu.pmem[3609] ;
wire \u_lsu.pmem[3610] ;
wire \u_lsu.pmem[3611] ;
wire \u_lsu.pmem[3612] ;
wire \u_lsu.pmem[3613] ;
wire \u_lsu.pmem[3614] ;
wire \u_lsu.pmem[3615] ;
wire \u_lsu.pmem[3616] ;
wire \u_lsu.pmem[3617] ;
wire \u_lsu.pmem[3618] ;
wire \u_lsu.pmem[3619] ;
wire \u_lsu.pmem[3620] ;
wire \u_lsu.pmem[3621] ;
wire \u_lsu.pmem[3622] ;
wire \u_lsu.pmem[3623] ;
wire \u_lsu.pmem[3624] ;
wire \u_lsu.pmem[3625] ;
wire \u_lsu.pmem[3626] ;
wire \u_lsu.pmem[3627] ;
wire \u_lsu.pmem[3628] ;
wire \u_lsu.pmem[3629] ;
wire \u_lsu.pmem[3630] ;
wire \u_lsu.pmem[3631] ;
wire \u_lsu.pmem[3632] ;
wire \u_lsu.pmem[3633] ;
wire \u_lsu.pmem[3634] ;
wire \u_lsu.pmem[3635] ;
wire \u_lsu.pmem[3636] ;
wire \u_lsu.pmem[3637] ;
wire \u_lsu.pmem[3638] ;
wire \u_lsu.pmem[3639] ;
wire \u_lsu.pmem[3640] ;
wire \u_lsu.pmem[3641] ;
wire \u_lsu.pmem[3642] ;
wire \u_lsu.pmem[3643] ;
wire \u_lsu.pmem[3644] ;
wire \u_lsu.pmem[3645] ;
wire \u_lsu.pmem[3646] ;
wire \u_lsu.pmem[3647] ;
wire \u_lsu.pmem[3648] ;
wire \u_lsu.pmem[3649] ;
wire \u_lsu.pmem[3650] ;
wire \u_lsu.pmem[3651] ;
wire \u_lsu.pmem[3652] ;
wire \u_lsu.pmem[3653] ;
wire \u_lsu.pmem[3654] ;
wire \u_lsu.pmem[3655] ;
wire \u_lsu.pmem[3656] ;
wire \u_lsu.pmem[3657] ;
wire \u_lsu.pmem[3658] ;
wire \u_lsu.pmem[3659] ;
wire \u_lsu.pmem[3660] ;
wire \u_lsu.pmem[3661] ;
wire \u_lsu.pmem[3662] ;
wire \u_lsu.pmem[3663] ;
wire \u_lsu.pmem[3664] ;
wire \u_lsu.pmem[3665] ;
wire \u_lsu.pmem[3666] ;
wire \u_lsu.pmem[3667] ;
wire \u_lsu.pmem[3668] ;
wire \u_lsu.pmem[3669] ;
wire \u_lsu.pmem[3670] ;
wire \u_lsu.pmem[3671] ;
wire \u_lsu.pmem[3672] ;
wire \u_lsu.pmem[3673] ;
wire \u_lsu.pmem[3674] ;
wire \u_lsu.pmem[3675] ;
wire \u_lsu.pmem[3676] ;
wire \u_lsu.pmem[3677] ;
wire \u_lsu.pmem[3678] ;
wire \u_lsu.pmem[3679] ;
wire \u_lsu.pmem[3680] ;
wire \u_lsu.pmem[3681] ;
wire \u_lsu.pmem[3682] ;
wire \u_lsu.pmem[3683] ;
wire \u_lsu.pmem[3684] ;
wire \u_lsu.pmem[3685] ;
wire \u_lsu.pmem[3686] ;
wire \u_lsu.pmem[3687] ;
wire \u_lsu.pmem[3688] ;
wire \u_lsu.pmem[3689] ;
wire \u_lsu.pmem[3690] ;
wire \u_lsu.pmem[3691] ;
wire \u_lsu.pmem[3692] ;
wire \u_lsu.pmem[3693] ;
wire \u_lsu.pmem[3694] ;
wire \u_lsu.pmem[3695] ;
wire \u_lsu.pmem[3696] ;
wire \u_lsu.pmem[3697] ;
wire \u_lsu.pmem[3698] ;
wire \u_lsu.pmem[3699] ;
wire \u_lsu.pmem[3700] ;
wire \u_lsu.pmem[3701] ;
wire \u_lsu.pmem[3702] ;
wire \u_lsu.pmem[3703] ;
wire \u_lsu.pmem[3704] ;
wire \u_lsu.pmem[3705] ;
wire \u_lsu.pmem[3706] ;
wire \u_lsu.pmem[3707] ;
wire \u_lsu.pmem[3708] ;
wire \u_lsu.pmem[3709] ;
wire \u_lsu.pmem[3710] ;
wire \u_lsu.pmem[3711] ;
wire \u_lsu.pmem[3712] ;
wire \u_lsu.pmem[3713] ;
wire \u_lsu.pmem[3714] ;
wire \u_lsu.pmem[3715] ;
wire \u_lsu.pmem[3716] ;
wire \u_lsu.pmem[3717] ;
wire \u_lsu.pmem[3718] ;
wire \u_lsu.pmem[3719] ;
wire \u_lsu.pmem[3720] ;
wire \u_lsu.pmem[3721] ;
wire \u_lsu.pmem[3722] ;
wire \u_lsu.pmem[3723] ;
wire \u_lsu.pmem[3724] ;
wire \u_lsu.pmem[3725] ;
wire \u_lsu.pmem[3726] ;
wire \u_lsu.pmem[3727] ;
wire \u_lsu.pmem[3728] ;
wire \u_lsu.pmem[3729] ;
wire \u_lsu.pmem[3730] ;
wire \u_lsu.pmem[3731] ;
wire \u_lsu.pmem[3732] ;
wire \u_lsu.pmem[3733] ;
wire \u_lsu.pmem[3734] ;
wire \u_lsu.pmem[3735] ;
wire \u_lsu.pmem[3736] ;
wire \u_lsu.pmem[3737] ;
wire \u_lsu.pmem[3738] ;
wire \u_lsu.pmem[3739] ;
wire \u_lsu.pmem[3740] ;
wire \u_lsu.pmem[3741] ;
wire \u_lsu.pmem[3742] ;
wire \u_lsu.pmem[3743] ;
wire \u_lsu.pmem[3744] ;
wire \u_lsu.pmem[3745] ;
wire \u_lsu.pmem[3746] ;
wire \u_lsu.pmem[3747] ;
wire \u_lsu.pmem[3748] ;
wire \u_lsu.pmem[3749] ;
wire \u_lsu.pmem[3750] ;
wire \u_lsu.pmem[3751] ;
wire \u_lsu.pmem[3752] ;
wire \u_lsu.pmem[3753] ;
wire \u_lsu.pmem[3754] ;
wire \u_lsu.pmem[3755] ;
wire \u_lsu.pmem[3756] ;
wire \u_lsu.pmem[3757] ;
wire \u_lsu.pmem[3758] ;
wire \u_lsu.pmem[3759] ;
wire \u_lsu.pmem[3760] ;
wire \u_lsu.pmem[3761] ;
wire \u_lsu.pmem[3762] ;
wire \u_lsu.pmem[3763] ;
wire \u_lsu.pmem[3764] ;
wire \u_lsu.pmem[3765] ;
wire \u_lsu.pmem[3766] ;
wire \u_lsu.pmem[3767] ;
wire \u_lsu.pmem[3768] ;
wire \u_lsu.pmem[3769] ;
wire \u_lsu.pmem[3770] ;
wire \u_lsu.pmem[3771] ;
wire \u_lsu.pmem[3772] ;
wire \u_lsu.pmem[3773] ;
wire \u_lsu.pmem[3774] ;
wire \u_lsu.pmem[3775] ;
wire \u_lsu.pmem[3776] ;
wire \u_lsu.pmem[3777] ;
wire \u_lsu.pmem[3778] ;
wire \u_lsu.pmem[3779] ;
wire \u_lsu.pmem[3780] ;
wire \u_lsu.pmem[3781] ;
wire \u_lsu.pmem[3782] ;
wire \u_lsu.pmem[3783] ;
wire \u_lsu.pmem[3784] ;
wire \u_lsu.pmem[3785] ;
wire \u_lsu.pmem[3786] ;
wire \u_lsu.pmem[3787] ;
wire \u_lsu.pmem[3788] ;
wire \u_lsu.pmem[3789] ;
wire \u_lsu.pmem[3790] ;
wire \u_lsu.pmem[3791] ;
wire \u_lsu.pmem[3792] ;
wire \u_lsu.pmem[3793] ;
wire \u_lsu.pmem[3794] ;
wire \u_lsu.pmem[3795] ;
wire \u_lsu.pmem[3796] ;
wire \u_lsu.pmem[3797] ;
wire \u_lsu.pmem[3798] ;
wire \u_lsu.pmem[3799] ;
wire \u_lsu.pmem[3800] ;
wire \u_lsu.pmem[3801] ;
wire \u_lsu.pmem[3802] ;
wire \u_lsu.pmem[3803] ;
wire \u_lsu.pmem[3804] ;
wire \u_lsu.pmem[3805] ;
wire \u_lsu.pmem[3806] ;
wire \u_lsu.pmem[3807] ;
wire \u_lsu.pmem[3808] ;
wire \u_lsu.pmem[3809] ;
wire \u_lsu.pmem[3810] ;
wire \u_lsu.pmem[3811] ;
wire \u_lsu.pmem[3812] ;
wire \u_lsu.pmem[3813] ;
wire \u_lsu.pmem[3814] ;
wire \u_lsu.pmem[3815] ;
wire \u_lsu.pmem[3816] ;
wire \u_lsu.pmem[3817] ;
wire \u_lsu.pmem[3818] ;
wire \u_lsu.pmem[3819] ;
wire \u_lsu.pmem[3820] ;
wire \u_lsu.pmem[3821] ;
wire \u_lsu.pmem[3822] ;
wire \u_lsu.pmem[3823] ;
wire \u_lsu.pmem[3824] ;
wire \u_lsu.pmem[3825] ;
wire \u_lsu.pmem[3826] ;
wire \u_lsu.pmem[3827] ;
wire \u_lsu.pmem[3828] ;
wire \u_lsu.pmem[3829] ;
wire \u_lsu.pmem[3830] ;
wire \u_lsu.pmem[3831] ;
wire \u_lsu.pmem[3832] ;
wire \u_lsu.pmem[3833] ;
wire \u_lsu.pmem[3834] ;
wire \u_lsu.pmem[3835] ;
wire \u_lsu.pmem[3836] ;
wire \u_lsu.pmem[3837] ;
wire \u_lsu.pmem[3838] ;
wire \u_lsu.pmem[3839] ;
wire \u_lsu.pmem[3840] ;
wire \u_lsu.pmem[3841] ;
wire \u_lsu.pmem[3842] ;
wire \u_lsu.pmem[3843] ;
wire \u_lsu.pmem[3844] ;
wire \u_lsu.pmem[3845] ;
wire \u_lsu.pmem[3846] ;
wire \u_lsu.pmem[3847] ;
wire \u_lsu.pmem[3848] ;
wire \u_lsu.pmem[3849] ;
wire \u_lsu.pmem[3850] ;
wire \u_lsu.pmem[3851] ;
wire \u_lsu.pmem[3852] ;
wire \u_lsu.pmem[3853] ;
wire \u_lsu.pmem[3854] ;
wire \u_lsu.pmem[3855] ;
wire \u_lsu.pmem[3856] ;
wire \u_lsu.pmem[3857] ;
wire \u_lsu.pmem[3858] ;
wire \u_lsu.pmem[3859] ;
wire \u_lsu.pmem[3860] ;
wire \u_lsu.pmem[3861] ;
wire \u_lsu.pmem[3862] ;
wire \u_lsu.pmem[3863] ;
wire \u_lsu.pmem[3864] ;
wire \u_lsu.pmem[3865] ;
wire \u_lsu.pmem[3866] ;
wire \u_lsu.pmem[3867] ;
wire \u_lsu.pmem[3868] ;
wire \u_lsu.pmem[3869] ;
wire \u_lsu.pmem[3870] ;
wire \u_lsu.pmem[3871] ;
wire \u_lsu.pmem[3872] ;
wire \u_lsu.pmem[3873] ;
wire \u_lsu.pmem[3874] ;
wire \u_lsu.pmem[3875] ;
wire \u_lsu.pmem[3876] ;
wire \u_lsu.pmem[3877] ;
wire \u_lsu.pmem[3878] ;
wire \u_lsu.pmem[3879] ;
wire \u_lsu.pmem[3880] ;
wire \u_lsu.pmem[3881] ;
wire \u_lsu.pmem[3882] ;
wire \u_lsu.pmem[3883] ;
wire \u_lsu.pmem[3884] ;
wire \u_lsu.pmem[3885] ;
wire \u_lsu.pmem[3886] ;
wire \u_lsu.pmem[3887] ;
wire \u_lsu.pmem[3888] ;
wire \u_lsu.pmem[3889] ;
wire \u_lsu.pmem[3890] ;
wire \u_lsu.pmem[3891] ;
wire \u_lsu.pmem[3892] ;
wire \u_lsu.pmem[3893] ;
wire \u_lsu.pmem[3894] ;
wire \u_lsu.pmem[3895] ;
wire \u_lsu.pmem[3896] ;
wire \u_lsu.pmem[3897] ;
wire \u_lsu.pmem[3898] ;
wire \u_lsu.pmem[3899] ;
wire \u_lsu.pmem[3900] ;
wire \u_lsu.pmem[3901] ;
wire \u_lsu.pmem[3902] ;
wire \u_lsu.pmem[3903] ;
wire \u_lsu.pmem[3904] ;
wire \u_lsu.pmem[3905] ;
wire \u_lsu.pmem[3906] ;
wire \u_lsu.pmem[3907] ;
wire \u_lsu.pmem[3908] ;
wire \u_lsu.pmem[3909] ;
wire \u_lsu.pmem[3910] ;
wire \u_lsu.pmem[3911] ;
wire \u_lsu.pmem[3912] ;
wire \u_lsu.pmem[3913] ;
wire \u_lsu.pmem[3914] ;
wire \u_lsu.pmem[3915] ;
wire \u_lsu.pmem[3916] ;
wire \u_lsu.pmem[3917] ;
wire \u_lsu.pmem[3918] ;
wire \u_lsu.pmem[3919] ;
wire \u_lsu.pmem[3920] ;
wire \u_lsu.pmem[3921] ;
wire \u_lsu.pmem[3922] ;
wire \u_lsu.pmem[3923] ;
wire \u_lsu.pmem[3924] ;
wire \u_lsu.pmem[3925] ;
wire \u_lsu.pmem[3926] ;
wire \u_lsu.pmem[3927] ;
wire \u_lsu.pmem[3928] ;
wire \u_lsu.pmem[3929] ;
wire \u_lsu.pmem[3930] ;
wire \u_lsu.pmem[3931] ;
wire \u_lsu.pmem[3932] ;
wire \u_lsu.pmem[3933] ;
wire \u_lsu.pmem[3934] ;
wire \u_lsu.pmem[3935] ;
wire \u_lsu.pmem[3936] ;
wire \u_lsu.pmem[3937] ;
wire \u_lsu.pmem[3938] ;
wire \u_lsu.pmem[3939] ;
wire \u_lsu.pmem[3940] ;
wire \u_lsu.pmem[3941] ;
wire \u_lsu.pmem[3942] ;
wire \u_lsu.pmem[3943] ;
wire \u_lsu.pmem[3944] ;
wire \u_lsu.pmem[3945] ;
wire \u_lsu.pmem[3946] ;
wire \u_lsu.pmem[3947] ;
wire \u_lsu.pmem[3948] ;
wire \u_lsu.pmem[3949] ;
wire \u_lsu.pmem[3950] ;
wire \u_lsu.pmem[3951] ;
wire \u_lsu.pmem[3952] ;
wire \u_lsu.pmem[3953] ;
wire \u_lsu.pmem[3954] ;
wire \u_lsu.pmem[3955] ;
wire \u_lsu.pmem[3956] ;
wire \u_lsu.pmem[3957] ;
wire \u_lsu.pmem[3958] ;
wire \u_lsu.pmem[3959] ;
wire \u_lsu.pmem[3960] ;
wire \u_lsu.pmem[3961] ;
wire \u_lsu.pmem[3962] ;
wire \u_lsu.pmem[3963] ;
wire \u_lsu.pmem[3964] ;
wire \u_lsu.pmem[3965] ;
wire \u_lsu.pmem[3966] ;
wire \u_lsu.pmem[3967] ;
wire \u_lsu.pmem[3968] ;
wire \u_lsu.pmem[3969] ;
wire \u_lsu.pmem[3970] ;
wire \u_lsu.pmem[3971] ;
wire \u_lsu.pmem[3972] ;
wire \u_lsu.pmem[3973] ;
wire \u_lsu.pmem[3974] ;
wire \u_lsu.pmem[3975] ;
wire \u_lsu.pmem[3976] ;
wire \u_lsu.pmem[3977] ;
wire \u_lsu.pmem[3978] ;
wire \u_lsu.pmem[3979] ;
wire \u_lsu.pmem[3980] ;
wire \u_lsu.pmem[3981] ;
wire \u_lsu.pmem[3982] ;
wire \u_lsu.pmem[3983] ;
wire \u_lsu.pmem[3984] ;
wire \u_lsu.pmem[3985] ;
wire \u_lsu.pmem[3986] ;
wire \u_lsu.pmem[3987] ;
wire \u_lsu.pmem[3988] ;
wire \u_lsu.pmem[3989] ;
wire \u_lsu.pmem[3990] ;
wire \u_lsu.pmem[3991] ;
wire \u_lsu.pmem[3992] ;
wire \u_lsu.pmem[3993] ;
wire \u_lsu.pmem[3994] ;
wire \u_lsu.pmem[3995] ;
wire \u_lsu.pmem[3996] ;
wire \u_lsu.pmem[3997] ;
wire \u_lsu.pmem[3998] ;
wire \u_lsu.pmem[3999] ;
wire \u_lsu.pmem[4000] ;
wire \u_lsu.pmem[4001] ;
wire \u_lsu.pmem[4002] ;
wire \u_lsu.pmem[4003] ;
wire \u_lsu.pmem[4004] ;
wire \u_lsu.pmem[4005] ;
wire \u_lsu.pmem[4006] ;
wire \u_lsu.pmem[4007] ;
wire \u_lsu.pmem[4008] ;
wire \u_lsu.pmem[4009] ;
wire \u_lsu.pmem[4010] ;
wire \u_lsu.pmem[4011] ;
wire \u_lsu.pmem[4012] ;
wire \u_lsu.pmem[4013] ;
wire \u_lsu.pmem[4014] ;
wire \u_lsu.pmem[4015] ;
wire \u_lsu.pmem[4016] ;
wire \u_lsu.pmem[4017] ;
wire \u_lsu.pmem[4018] ;
wire \u_lsu.pmem[4019] ;
wire \u_lsu.pmem[4020] ;
wire \u_lsu.pmem[4021] ;
wire \u_lsu.pmem[4022] ;
wire \u_lsu.pmem[4023] ;
wire \u_lsu.pmem[4024] ;
wire \u_lsu.pmem[4025] ;
wire \u_lsu.pmem[4026] ;
wire \u_lsu.pmem[4027] ;
wire \u_lsu.pmem[4028] ;
wire \u_lsu.pmem[4029] ;
wire \u_lsu.pmem[4030] ;
wire \u_lsu.pmem[4031] ;
wire \u_lsu.pmem[4032] ;
wire \u_lsu.pmem[4033] ;
wire \u_lsu.pmem[4034] ;
wire \u_lsu.pmem[4035] ;
wire \u_lsu.pmem[4036] ;
wire \u_lsu.pmem[4037] ;
wire \u_lsu.pmem[4038] ;
wire \u_lsu.pmem[4039] ;
wire \u_lsu.pmem[4040] ;
wire \u_lsu.pmem[4041] ;
wire \u_lsu.pmem[4042] ;
wire \u_lsu.pmem[4043] ;
wire \u_lsu.pmem[4044] ;
wire \u_lsu.pmem[4045] ;
wire \u_lsu.pmem[4046] ;
wire \u_lsu.pmem[4047] ;
wire \u_lsu.pmem[4048] ;
wire \u_lsu.pmem[4049] ;
wire \u_lsu.pmem[4050] ;
wire \u_lsu.pmem[4051] ;
wire \u_lsu.pmem[4052] ;
wire \u_lsu.pmem[4053] ;
wire \u_lsu.pmem[4054] ;
wire \u_lsu.pmem[4055] ;
wire \u_lsu.pmem[4056] ;
wire \u_lsu.pmem[4057] ;
wire \u_lsu.pmem[4058] ;
wire \u_lsu.pmem[4059] ;
wire \u_lsu.pmem[4060] ;
wire \u_lsu.pmem[4061] ;
wire \u_lsu.pmem[4062] ;
wire \u_lsu.pmem[4063] ;
wire \u_lsu.pmem[4064] ;
wire \u_lsu.pmem[4065] ;
wire \u_lsu.pmem[4066] ;
wire \u_lsu.pmem[4067] ;
wire \u_lsu.pmem[4068] ;
wire \u_lsu.pmem[4069] ;
wire \u_lsu.pmem[4070] ;
wire \u_lsu.pmem[4071] ;
wire \u_lsu.pmem[4072] ;
wire \u_lsu.pmem[4073] ;
wire \u_lsu.pmem[4074] ;
wire \u_lsu.pmem[4075] ;
wire \u_lsu.pmem[4076] ;
wire \u_lsu.pmem[4077] ;
wire \u_lsu.pmem[4078] ;
wire \u_lsu.pmem[4079] ;
wire \u_lsu.pmem[4080] ;
wire \u_lsu.pmem[4081] ;
wire \u_lsu.pmem[4082] ;
wire \u_lsu.pmem[4083] ;
wire \u_lsu.pmem[4084] ;
wire \u_lsu.pmem[4085] ;
wire \u_lsu.pmem[4086] ;
wire \u_lsu.pmem[4087] ;
wire \u_lsu.pmem[4088] ;
wire \u_lsu.pmem[4089] ;
wire \u_lsu.pmem[4090] ;
wire \u_lsu.pmem[4091] ;
wire \u_lsu.pmem[4092] ;
wire \u_lsu.pmem[4093] ;
wire \u_lsu.pmem[4094] ;
wire \u_lsu.pmem[4095] ;
wire \u_lsu.pmem[4096] ;
wire \u_lsu.pmem[4097] ;
wire \u_lsu.pmem[4098] ;
wire \u_lsu.pmem[4099] ;
wire \u_lsu.pmem[4100] ;
wire \u_lsu.pmem[4101] ;
wire \u_lsu.pmem[4102] ;
wire \u_lsu.pmem[4103] ;
wire \u_lsu.pmem[4104] ;
wire \u_lsu.pmem[4105] ;
wire \u_lsu.pmem[4106] ;
wire \u_lsu.pmem[4107] ;
wire \u_lsu.pmem[4108] ;
wire \u_lsu.pmem[4109] ;
wire \u_lsu.pmem[4110] ;
wire \u_lsu.pmem[4111] ;
wire \u_lsu.pmem[4112] ;
wire \u_lsu.pmem[4113] ;
wire \u_lsu.pmem[4114] ;
wire \u_lsu.pmem[4115] ;
wire \u_lsu.pmem[4116] ;
wire \u_lsu.pmem[4117] ;
wire \u_lsu.pmem[4118] ;
wire \u_lsu.pmem[4119] ;
wire \u_lsu.pmem[4120] ;
wire \u_lsu.pmem[4121] ;
wire \u_lsu.pmem[4122] ;
wire \u_lsu.pmem[4123] ;
wire \u_lsu.pmem[4124] ;
wire \u_lsu.pmem[4125] ;
wire \u_lsu.pmem[4126] ;
wire \u_lsu.pmem[4127] ;
wire \u_lsu.pmem[4128] ;
wire \u_lsu.pmem[4129] ;
wire \u_lsu.pmem[4130] ;
wire \u_lsu.pmem[4131] ;
wire \u_lsu.pmem[4132] ;
wire \u_lsu.pmem[4133] ;
wire \u_lsu.pmem[4134] ;
wire \u_lsu.pmem[4135] ;
wire \u_lsu.pmem[4136] ;
wire \u_lsu.pmem[4137] ;
wire \u_lsu.pmem[4138] ;
wire \u_lsu.pmem[4139] ;
wire \u_lsu.pmem[4140] ;
wire \u_lsu.pmem[4141] ;
wire \u_lsu.pmem[4142] ;
wire \u_lsu.pmem[4143] ;
wire \u_lsu.pmem[4144] ;
wire \u_lsu.pmem[4145] ;
wire \u_lsu.pmem[4146] ;
wire \u_lsu.pmem[4147] ;
wire \u_lsu.pmem[4148] ;
wire \u_lsu.pmem[4149] ;
wire \u_lsu.pmem[4150] ;
wire \u_lsu.pmem[4151] ;
wire \u_lsu.pmem[4152] ;
wire \u_lsu.pmem[4153] ;
wire \u_lsu.pmem[4154] ;
wire \u_lsu.pmem[4155] ;
wire \u_lsu.pmem[4156] ;
wire \u_lsu.pmem[4157] ;
wire \u_lsu.pmem[4158] ;
wire \u_lsu.pmem[4159] ;
wire \u_lsu.pmem[4160] ;
wire \u_lsu.pmem[4161] ;
wire \u_lsu.pmem[4162] ;
wire \u_lsu.pmem[4163] ;
wire \u_lsu.pmem[4164] ;
wire \u_lsu.pmem[4165] ;
wire \u_lsu.pmem[4166] ;
wire \u_lsu.pmem[4167] ;
wire \u_lsu.pmem[4168] ;
wire \u_lsu.pmem[4169] ;
wire \u_lsu.pmem[4170] ;
wire \u_lsu.pmem[4171] ;
wire \u_lsu.pmem[4172] ;
wire \u_lsu.pmem[4173] ;
wire \u_lsu.pmem[4174] ;
wire \u_lsu.pmem[4175] ;
wire \u_lsu.pmem[4176] ;
wire \u_lsu.pmem[4177] ;
wire \u_lsu.pmem[4178] ;
wire \u_lsu.pmem[4179] ;
wire \u_lsu.pmem[4180] ;
wire \u_lsu.pmem[4181] ;
wire \u_lsu.pmem[4182] ;
wire \u_lsu.pmem[4183] ;
wire \u_lsu.pmem[4184] ;
wire \u_lsu.pmem[4185] ;
wire \u_lsu.pmem[4186] ;
wire \u_lsu.pmem[4187] ;
wire \u_lsu.pmem[4188] ;
wire \u_lsu.pmem[4189] ;
wire \u_lsu.pmem[4190] ;
wire \u_lsu.pmem[4191] ;
wire \u_lsu.pmem[4192] ;
wire \u_lsu.pmem[4193] ;
wire \u_lsu.pmem[4194] ;
wire \u_lsu.pmem[4195] ;
wire \u_lsu.pmem[4196] ;
wire \u_lsu.pmem[4197] ;
wire \u_lsu.pmem[4198] ;
wire \u_lsu.pmem[4199] ;
wire \u_lsu.pmem[4200] ;
wire \u_lsu.pmem[4201] ;
wire \u_lsu.pmem[4202] ;
wire \u_lsu.pmem[4203] ;
wire \u_lsu.pmem[4204] ;
wire \u_lsu.pmem[4205] ;
wire \u_lsu.pmem[4206] ;
wire \u_lsu.pmem[4207] ;
wire \u_lsu.pmem[4208] ;
wire \u_lsu.pmem[4209] ;
wire \u_lsu.pmem[4210] ;
wire \u_lsu.pmem[4211] ;
wire \u_lsu.pmem[4212] ;
wire \u_lsu.pmem[4213] ;
wire \u_lsu.pmem[4214] ;
wire \u_lsu.pmem[4215] ;
wire \u_lsu.pmem[4216] ;
wire \u_lsu.pmem[4217] ;
wire \u_lsu.pmem[4218] ;
wire \u_lsu.pmem[4219] ;
wire \u_lsu.pmem[4220] ;
wire \u_lsu.pmem[4221] ;
wire \u_lsu.pmem[4222] ;
wire \u_lsu.pmem[4223] ;
wire \u_lsu.pmem[4224] ;
wire \u_lsu.pmem[4225] ;
wire \u_lsu.pmem[4226] ;
wire \u_lsu.pmem[4227] ;
wire \u_lsu.pmem[4228] ;
wire \u_lsu.pmem[4229] ;
wire \u_lsu.pmem[4230] ;
wire \u_lsu.pmem[4231] ;
wire \u_lsu.pmem[4232] ;
wire \u_lsu.pmem[4233] ;
wire \u_lsu.pmem[4234] ;
wire \u_lsu.pmem[4235] ;
wire \u_lsu.pmem[4236] ;
wire \u_lsu.pmem[4237] ;
wire \u_lsu.pmem[4238] ;
wire \u_lsu.pmem[4239] ;
wire \u_lsu.pmem[4240] ;
wire \u_lsu.pmem[4241] ;
wire \u_lsu.pmem[4242] ;
wire \u_lsu.pmem[4243] ;
wire \u_lsu.pmem[4244] ;
wire \u_lsu.pmem[4245] ;
wire \u_lsu.pmem[4246] ;
wire \u_lsu.pmem[4247] ;
wire \u_lsu.pmem[4248] ;
wire \u_lsu.pmem[4249] ;
wire \u_lsu.pmem[4250] ;
wire \u_lsu.pmem[4251] ;
wire \u_lsu.pmem[4252] ;
wire \u_lsu.pmem[4253] ;
wire \u_lsu.pmem[4254] ;
wire \u_lsu.pmem[4255] ;
wire \u_lsu.pmem[4256] ;
wire \u_lsu.pmem[4257] ;
wire \u_lsu.pmem[4258] ;
wire \u_lsu.pmem[4259] ;
wire \u_lsu.pmem[4260] ;
wire \u_lsu.pmem[4261] ;
wire \u_lsu.pmem[4262] ;
wire \u_lsu.pmem[4263] ;
wire \u_lsu.pmem[4264] ;
wire \u_lsu.pmem[4265] ;
wire \u_lsu.pmem[4266] ;
wire \u_lsu.pmem[4267] ;
wire \u_lsu.pmem[4268] ;
wire \u_lsu.pmem[4269] ;
wire \u_lsu.pmem[4270] ;
wire \u_lsu.pmem[4271] ;
wire \u_lsu.pmem[4272] ;
wire \u_lsu.pmem[4273] ;
wire \u_lsu.pmem[4274] ;
wire \u_lsu.pmem[4275] ;
wire \u_lsu.pmem[4276] ;
wire \u_lsu.pmem[4277] ;
wire \u_lsu.pmem[4278] ;
wire \u_lsu.pmem[4279] ;
wire \u_lsu.pmem[4280] ;
wire \u_lsu.pmem[4281] ;
wire \u_lsu.pmem[4282] ;
wire \u_lsu.pmem[4283] ;
wire \u_lsu.pmem[4284] ;
wire \u_lsu.pmem[4285] ;
wire \u_lsu.pmem[4286] ;
wire \u_lsu.pmem[4287] ;
wire \u_lsu.pmem[4288] ;
wire \u_lsu.pmem[4289] ;
wire \u_lsu.pmem[4290] ;
wire \u_lsu.pmem[4291] ;
wire \u_lsu.pmem[4292] ;
wire \u_lsu.pmem[4293] ;
wire \u_lsu.pmem[4294] ;
wire \u_lsu.pmem[4295] ;
wire \u_lsu.pmem[4296] ;
wire \u_lsu.pmem[4297] ;
wire \u_lsu.pmem[4298] ;
wire \u_lsu.pmem[4299] ;
wire \u_lsu.pmem[4300] ;
wire \u_lsu.pmem[4301] ;
wire \u_lsu.pmem[4302] ;
wire \u_lsu.pmem[4303] ;
wire \u_lsu.pmem[4304] ;
wire \u_lsu.pmem[4305] ;
wire \u_lsu.pmem[4306] ;
wire \u_lsu.pmem[4307] ;
wire \u_lsu.pmem[4308] ;
wire \u_lsu.pmem[4309] ;
wire \u_lsu.pmem[4310] ;
wire \u_lsu.pmem[4311] ;
wire \u_lsu.pmem[4312] ;
wire \u_lsu.pmem[4313] ;
wire \u_lsu.pmem[4314] ;
wire \u_lsu.pmem[4315] ;
wire \u_lsu.pmem[4316] ;
wire \u_lsu.pmem[4317] ;
wire \u_lsu.pmem[4318] ;
wire \u_lsu.pmem[4319] ;
wire \u_lsu.pmem[4320] ;
wire \u_lsu.pmem[4321] ;
wire \u_lsu.pmem[4322] ;
wire \u_lsu.pmem[4323] ;
wire \u_lsu.pmem[4324] ;
wire \u_lsu.pmem[4325] ;
wire \u_lsu.pmem[4326] ;
wire \u_lsu.pmem[4327] ;
wire \u_lsu.pmem[4328] ;
wire \u_lsu.pmem[4329] ;
wire \u_lsu.pmem[4330] ;
wire \u_lsu.pmem[4331] ;
wire \u_lsu.pmem[4332] ;
wire \u_lsu.pmem[4333] ;
wire \u_lsu.pmem[4334] ;
wire \u_lsu.pmem[4335] ;
wire \u_lsu.pmem[4336] ;
wire \u_lsu.pmem[4337] ;
wire \u_lsu.pmem[4338] ;
wire \u_lsu.pmem[4339] ;
wire \u_lsu.pmem[4340] ;
wire \u_lsu.pmem[4341] ;
wire \u_lsu.pmem[4342] ;
wire \u_lsu.pmem[4343] ;
wire \u_lsu.pmem[4344] ;
wire \u_lsu.pmem[4345] ;
wire \u_lsu.pmem[4346] ;
wire \u_lsu.pmem[4347] ;
wire \u_lsu.pmem[4348] ;
wire \u_lsu.pmem[4349] ;
wire \u_lsu.pmem[4350] ;
wire \u_lsu.pmem[4351] ;
wire \u_lsu.pmem[4352] ;
wire \u_lsu.pmem[4353] ;
wire \u_lsu.pmem[4354] ;
wire \u_lsu.pmem[4355] ;
wire \u_lsu.pmem[4356] ;
wire \u_lsu.pmem[4357] ;
wire \u_lsu.pmem[4358] ;
wire \u_lsu.pmem[4359] ;
wire \u_lsu.pmem[4360] ;
wire \u_lsu.pmem[4361] ;
wire \u_lsu.pmem[4362] ;
wire \u_lsu.pmem[4363] ;
wire \u_lsu.pmem[4364] ;
wire \u_lsu.pmem[4365] ;
wire \u_lsu.pmem[4366] ;
wire \u_lsu.pmem[4367] ;
wire \u_lsu.pmem[4368] ;
wire \u_lsu.pmem[4369] ;
wire \u_lsu.pmem[4370] ;
wire \u_lsu.pmem[4371] ;
wire \u_lsu.pmem[4372] ;
wire \u_lsu.pmem[4373] ;
wire \u_lsu.pmem[4374] ;
wire \u_lsu.pmem[4375] ;
wire \u_lsu.pmem[4376] ;
wire \u_lsu.pmem[4377] ;
wire \u_lsu.pmem[4378] ;
wire \u_lsu.pmem[4379] ;
wire \u_lsu.pmem[4380] ;
wire \u_lsu.pmem[4381] ;
wire \u_lsu.pmem[4382] ;
wire \u_lsu.pmem[4383] ;
wire \u_lsu.pmem[4384] ;
wire \u_lsu.pmem[4385] ;
wire \u_lsu.pmem[4386] ;
wire \u_lsu.pmem[4387] ;
wire \u_lsu.pmem[4388] ;
wire \u_lsu.pmem[4389] ;
wire \u_lsu.pmem[4390] ;
wire \u_lsu.pmem[4391] ;
wire \u_lsu.pmem[4392] ;
wire \u_lsu.pmem[4393] ;
wire \u_lsu.pmem[4394] ;
wire \u_lsu.pmem[4395] ;
wire \u_lsu.pmem[4396] ;
wire \u_lsu.pmem[4397] ;
wire \u_lsu.pmem[4398] ;
wire \u_lsu.pmem[4399] ;
wire \u_lsu.pmem[4400] ;
wire \u_lsu.pmem[4401] ;
wire \u_lsu.pmem[4402] ;
wire \u_lsu.pmem[4403] ;
wire \u_lsu.pmem[4404] ;
wire \u_lsu.pmem[4405] ;
wire \u_lsu.pmem[4406] ;
wire \u_lsu.pmem[4407] ;
wire \u_lsu.pmem[4408] ;
wire \u_lsu.pmem[4409] ;
wire \u_lsu.pmem[4410] ;
wire \u_lsu.pmem[4411] ;
wire \u_lsu.pmem[4412] ;
wire \u_lsu.pmem[4413] ;
wire \u_lsu.pmem[4414] ;
wire \u_lsu.pmem[4415] ;
wire \u_lsu.pmem[4416] ;
wire \u_lsu.pmem[4417] ;
wire \u_lsu.pmem[4418] ;
wire \u_lsu.pmem[4419] ;
wire \u_lsu.pmem[4420] ;
wire \u_lsu.pmem[4421] ;
wire \u_lsu.pmem[4422] ;
wire \u_lsu.pmem[4423] ;
wire \u_lsu.pmem[4424] ;
wire \u_lsu.pmem[4425] ;
wire \u_lsu.pmem[4426] ;
wire \u_lsu.pmem[4427] ;
wire \u_lsu.pmem[4428] ;
wire \u_lsu.pmem[4429] ;
wire \u_lsu.pmem[4430] ;
wire \u_lsu.pmem[4431] ;
wire \u_lsu.pmem[4432] ;
wire \u_lsu.pmem[4433] ;
wire \u_lsu.pmem[4434] ;
wire \u_lsu.pmem[4435] ;
wire \u_lsu.pmem[4436] ;
wire \u_lsu.pmem[4437] ;
wire \u_lsu.pmem[4438] ;
wire \u_lsu.pmem[4439] ;
wire \u_lsu.pmem[4440] ;
wire \u_lsu.pmem[4441] ;
wire \u_lsu.pmem[4442] ;
wire \u_lsu.pmem[4443] ;
wire \u_lsu.pmem[4444] ;
wire \u_lsu.pmem[4445] ;
wire \u_lsu.pmem[4446] ;
wire \u_lsu.pmem[4447] ;
wire \u_lsu.pmem[4448] ;
wire \u_lsu.pmem[4449] ;
wire \u_lsu.pmem[4450] ;
wire \u_lsu.pmem[4451] ;
wire \u_lsu.pmem[4452] ;
wire \u_lsu.pmem[4453] ;
wire \u_lsu.pmem[4454] ;
wire \u_lsu.pmem[4455] ;
wire \u_lsu.pmem[4456] ;
wire \u_lsu.pmem[4457] ;
wire \u_lsu.pmem[4458] ;
wire \u_lsu.pmem[4459] ;
wire \u_lsu.pmem[4460] ;
wire \u_lsu.pmem[4461] ;
wire \u_lsu.pmem[4462] ;
wire \u_lsu.pmem[4463] ;
wire \u_lsu.pmem[4464] ;
wire \u_lsu.pmem[4465] ;
wire \u_lsu.pmem[4466] ;
wire \u_lsu.pmem[4467] ;
wire \u_lsu.pmem[4468] ;
wire \u_lsu.pmem[4469] ;
wire \u_lsu.pmem[4470] ;
wire \u_lsu.pmem[4471] ;
wire \u_lsu.pmem[4472] ;
wire \u_lsu.pmem[4473] ;
wire \u_lsu.pmem[4474] ;
wire \u_lsu.pmem[4475] ;
wire \u_lsu.pmem[4476] ;
wire \u_lsu.pmem[4477] ;
wire \u_lsu.pmem[4478] ;
wire \u_lsu.pmem[4479] ;
wire \u_lsu.pmem[4480] ;
wire \u_lsu.pmem[4481] ;
wire \u_lsu.pmem[4482] ;
wire \u_lsu.pmem[4483] ;
wire \u_lsu.pmem[4484] ;
wire \u_lsu.pmem[4485] ;
wire \u_lsu.pmem[4486] ;
wire \u_lsu.pmem[4487] ;
wire \u_lsu.pmem[4488] ;
wire \u_lsu.pmem[4489] ;
wire \u_lsu.pmem[4490] ;
wire \u_lsu.pmem[4491] ;
wire \u_lsu.pmem[4492] ;
wire \u_lsu.pmem[4493] ;
wire \u_lsu.pmem[4494] ;
wire \u_lsu.pmem[4495] ;
wire \u_lsu.pmem[4496] ;
wire \u_lsu.pmem[4497] ;
wire \u_lsu.pmem[4498] ;
wire \u_lsu.pmem[4499] ;
wire \u_lsu.pmem[4500] ;
wire \u_lsu.pmem[4501] ;
wire \u_lsu.pmem[4502] ;
wire \u_lsu.pmem[4503] ;
wire \u_lsu.pmem[4504] ;
wire \u_lsu.pmem[4505] ;
wire \u_lsu.pmem[4506] ;
wire \u_lsu.pmem[4507] ;
wire \u_lsu.pmem[4508] ;
wire \u_lsu.pmem[4509] ;
wire \u_lsu.pmem[4510] ;
wire \u_lsu.pmem[4511] ;
wire \u_lsu.pmem[4512] ;
wire \u_lsu.pmem[4513] ;
wire \u_lsu.pmem[4514] ;
wire \u_lsu.pmem[4515] ;
wire \u_lsu.pmem[4516] ;
wire \u_lsu.pmem[4517] ;
wire \u_lsu.pmem[4518] ;
wire \u_lsu.pmem[4519] ;
wire \u_lsu.pmem[4520] ;
wire \u_lsu.pmem[4521] ;
wire \u_lsu.pmem[4522] ;
wire \u_lsu.pmem[4523] ;
wire \u_lsu.pmem[4524] ;
wire \u_lsu.pmem[4525] ;
wire \u_lsu.pmem[4526] ;
wire \u_lsu.pmem[4527] ;
wire \u_lsu.pmem[4528] ;
wire \u_lsu.pmem[4529] ;
wire \u_lsu.pmem[4530] ;
wire \u_lsu.pmem[4531] ;
wire \u_lsu.pmem[4532] ;
wire \u_lsu.pmem[4533] ;
wire \u_lsu.pmem[4534] ;
wire \u_lsu.pmem[4535] ;
wire \u_lsu.pmem[4536] ;
wire \u_lsu.pmem[4537] ;
wire \u_lsu.pmem[4538] ;
wire \u_lsu.pmem[4539] ;
wire \u_lsu.pmem[4540] ;
wire \u_lsu.pmem[4541] ;
wire \u_lsu.pmem[4542] ;
wire \u_lsu.pmem[4543] ;
wire \u_lsu.pmem[4544] ;
wire \u_lsu.pmem[4545] ;
wire \u_lsu.pmem[4546] ;
wire \u_lsu.pmem[4547] ;
wire \u_lsu.pmem[4548] ;
wire \u_lsu.pmem[4549] ;
wire \u_lsu.pmem[4550] ;
wire \u_lsu.pmem[4551] ;
wire \u_lsu.pmem[4552] ;
wire \u_lsu.pmem[4553] ;
wire \u_lsu.pmem[4554] ;
wire \u_lsu.pmem[4555] ;
wire \u_lsu.pmem[4556] ;
wire \u_lsu.pmem[4557] ;
wire \u_lsu.pmem[4558] ;
wire \u_lsu.pmem[4559] ;
wire \u_lsu.pmem[4560] ;
wire \u_lsu.pmem[4561] ;
wire \u_lsu.pmem[4562] ;
wire \u_lsu.pmem[4563] ;
wire \u_lsu.pmem[4564] ;
wire \u_lsu.pmem[4565] ;
wire \u_lsu.pmem[4566] ;
wire \u_lsu.pmem[4567] ;
wire \u_lsu.pmem[4568] ;
wire \u_lsu.pmem[4569] ;
wire \u_lsu.pmem[4570] ;
wire \u_lsu.pmem[4571] ;
wire \u_lsu.pmem[4572] ;
wire \u_lsu.pmem[4573] ;
wire \u_lsu.pmem[4574] ;
wire \u_lsu.pmem[4575] ;
wire \u_lsu.pmem[4576] ;
wire \u_lsu.pmem[4577] ;
wire \u_lsu.pmem[4578] ;
wire \u_lsu.pmem[4579] ;
wire \u_lsu.pmem[4580] ;
wire \u_lsu.pmem[4581] ;
wire \u_lsu.pmem[4582] ;
wire \u_lsu.pmem[4583] ;
wire \u_lsu.pmem[4584] ;
wire \u_lsu.pmem[4585] ;
wire \u_lsu.pmem[4586] ;
wire \u_lsu.pmem[4587] ;
wire \u_lsu.pmem[4588] ;
wire \u_lsu.pmem[4589] ;
wire \u_lsu.pmem[4590] ;
wire \u_lsu.pmem[4591] ;
wire \u_lsu.pmem[4592] ;
wire \u_lsu.pmem[4593] ;
wire \u_lsu.pmem[4594] ;
wire \u_lsu.pmem[4595] ;
wire \u_lsu.pmem[4596] ;
wire \u_lsu.pmem[4597] ;
wire \u_lsu.pmem[4598] ;
wire \u_lsu.pmem[4599] ;
wire \u_lsu.pmem[4600] ;
wire \u_lsu.pmem[4601] ;
wire \u_lsu.pmem[4602] ;
wire \u_lsu.pmem[4603] ;
wire \u_lsu.pmem[4604] ;
wire \u_lsu.pmem[4605] ;
wire \u_lsu.pmem[4606] ;
wire \u_lsu.pmem[4607] ;
wire \u_lsu.pmem[4608] ;
wire \u_lsu.pmem[4609] ;
wire \u_lsu.pmem[4610] ;
wire \u_lsu.pmem[4611] ;
wire \u_lsu.pmem[4612] ;
wire \u_lsu.pmem[4613] ;
wire \u_lsu.pmem[4614] ;
wire \u_lsu.pmem[4615] ;
wire \u_lsu.pmem[4616] ;
wire \u_lsu.pmem[4617] ;
wire \u_lsu.pmem[4618] ;
wire \u_lsu.pmem[4619] ;
wire \u_lsu.pmem[4620] ;
wire \u_lsu.pmem[4621] ;
wire \u_lsu.pmem[4622] ;
wire \u_lsu.pmem[4623] ;
wire \u_lsu.pmem[4624] ;
wire \u_lsu.pmem[4625] ;
wire \u_lsu.pmem[4626] ;
wire \u_lsu.pmem[4627] ;
wire \u_lsu.pmem[4628] ;
wire \u_lsu.pmem[4629] ;
wire \u_lsu.pmem[4630] ;
wire \u_lsu.pmem[4631] ;
wire \u_lsu.pmem[4632] ;
wire \u_lsu.pmem[4633] ;
wire \u_lsu.pmem[4634] ;
wire \u_lsu.pmem[4635] ;
wire \u_lsu.pmem[4636] ;
wire \u_lsu.pmem[4637] ;
wire \u_lsu.pmem[4638] ;
wire \u_lsu.pmem[4639] ;
wire \u_lsu.pmem[4640] ;
wire \u_lsu.pmem[4641] ;
wire \u_lsu.pmem[4642] ;
wire \u_lsu.pmem[4643] ;
wire \u_lsu.pmem[4644] ;
wire \u_lsu.pmem[4645] ;
wire \u_lsu.pmem[4646] ;
wire \u_lsu.pmem[4647] ;
wire \u_lsu.pmem[4648] ;
wire \u_lsu.pmem[4649] ;
wire \u_lsu.pmem[4650] ;
wire \u_lsu.pmem[4651] ;
wire \u_lsu.pmem[4652] ;
wire \u_lsu.pmem[4653] ;
wire \u_lsu.pmem[4654] ;
wire \u_lsu.pmem[4655] ;
wire \u_lsu.pmem[4656] ;
wire \u_lsu.pmem[4657] ;
wire \u_lsu.pmem[4658] ;
wire \u_lsu.pmem[4659] ;
wire \u_lsu.pmem[4660] ;
wire \u_lsu.pmem[4661] ;
wire \u_lsu.pmem[4662] ;
wire \u_lsu.pmem[4663] ;
wire \u_lsu.pmem[4664] ;
wire \u_lsu.pmem[4665] ;
wire \u_lsu.pmem[4666] ;
wire \u_lsu.pmem[4667] ;
wire \u_lsu.pmem[4668] ;
wire \u_lsu.pmem[4669] ;
wire \u_lsu.pmem[4670] ;
wire \u_lsu.pmem[4671] ;
wire \u_lsu.pmem[4672] ;
wire \u_lsu.pmem[4673] ;
wire \u_lsu.pmem[4674] ;
wire \u_lsu.pmem[4675] ;
wire \u_lsu.pmem[4676] ;
wire \u_lsu.pmem[4677] ;
wire \u_lsu.pmem[4678] ;
wire \u_lsu.pmem[4679] ;
wire \u_lsu.pmem[4680] ;
wire \u_lsu.pmem[4681] ;
wire \u_lsu.pmem[4682] ;
wire \u_lsu.pmem[4683] ;
wire \u_lsu.pmem[4684] ;
wire \u_lsu.pmem[4685] ;
wire \u_lsu.pmem[4686] ;
wire \u_lsu.pmem[4687] ;
wire \u_lsu.pmem[4688] ;
wire \u_lsu.pmem[4689] ;
wire \u_lsu.pmem[4690] ;
wire \u_lsu.pmem[4691] ;
wire \u_lsu.pmem[4692] ;
wire \u_lsu.pmem[4693] ;
wire \u_lsu.pmem[4694] ;
wire \u_lsu.pmem[4695] ;
wire \u_lsu.pmem[4696] ;
wire \u_lsu.pmem[4697] ;
wire \u_lsu.pmem[4698] ;
wire \u_lsu.pmem[4699] ;
wire \u_lsu.pmem[4700] ;
wire \u_lsu.pmem[4701] ;
wire \u_lsu.pmem[4702] ;
wire \u_lsu.pmem[4703] ;
wire \u_lsu.pmem[4704] ;
wire \u_lsu.pmem[4705] ;
wire \u_lsu.pmem[4706] ;
wire \u_lsu.pmem[4707] ;
wire \u_lsu.pmem[4708] ;
wire \u_lsu.pmem[4709] ;
wire \u_lsu.pmem[4710] ;
wire \u_lsu.pmem[4711] ;
wire \u_lsu.pmem[4712] ;
wire \u_lsu.pmem[4713] ;
wire \u_lsu.pmem[4714] ;
wire \u_lsu.pmem[4715] ;
wire \u_lsu.pmem[4716] ;
wire \u_lsu.pmem[4717] ;
wire \u_lsu.pmem[4718] ;
wire \u_lsu.pmem[4719] ;
wire \u_lsu.pmem[4720] ;
wire \u_lsu.pmem[4721] ;
wire \u_lsu.pmem[4722] ;
wire \u_lsu.pmem[4723] ;
wire \u_lsu.pmem[4724] ;
wire \u_lsu.pmem[4725] ;
wire \u_lsu.pmem[4726] ;
wire \u_lsu.pmem[4727] ;
wire \u_lsu.pmem[4728] ;
wire \u_lsu.pmem[4729] ;
wire \u_lsu.pmem[4730] ;
wire \u_lsu.pmem[4731] ;
wire \u_lsu.pmem[4732] ;
wire \u_lsu.pmem[4733] ;
wire \u_lsu.pmem[4734] ;
wire \u_lsu.pmem[4735] ;
wire \u_lsu.pmem[4736] ;
wire \u_lsu.pmem[4737] ;
wire \u_lsu.pmem[4738] ;
wire \u_lsu.pmem[4739] ;
wire \u_lsu.pmem[4740] ;
wire \u_lsu.pmem[4741] ;
wire \u_lsu.pmem[4742] ;
wire \u_lsu.pmem[4743] ;
wire \u_lsu.pmem[4744] ;
wire \u_lsu.pmem[4745] ;
wire \u_lsu.pmem[4746] ;
wire \u_lsu.pmem[4747] ;
wire \u_lsu.pmem[4748] ;
wire \u_lsu.pmem[4749] ;
wire \u_lsu.pmem[4750] ;
wire \u_lsu.pmem[4751] ;
wire \u_lsu.pmem[4752] ;
wire \u_lsu.pmem[4753] ;
wire \u_lsu.pmem[4754] ;
wire \u_lsu.pmem[4755] ;
wire \u_lsu.pmem[4756] ;
wire \u_lsu.pmem[4757] ;
wire \u_lsu.pmem[4758] ;
wire \u_lsu.pmem[4759] ;
wire \u_lsu.pmem[4760] ;
wire \u_lsu.pmem[4761] ;
wire \u_lsu.pmem[4762] ;
wire \u_lsu.pmem[4763] ;
wire \u_lsu.pmem[4764] ;
wire \u_lsu.pmem[4765] ;
wire \u_lsu.pmem[4766] ;
wire \u_lsu.pmem[4767] ;
wire \u_lsu.pmem[4768] ;
wire \u_lsu.pmem[4769] ;
wire \u_lsu.pmem[4770] ;
wire \u_lsu.pmem[4771] ;
wire \u_lsu.pmem[4772] ;
wire \u_lsu.pmem[4773] ;
wire \u_lsu.pmem[4774] ;
wire \u_lsu.pmem[4775] ;
wire \u_lsu.pmem[4776] ;
wire \u_lsu.pmem[4777] ;
wire \u_lsu.pmem[4778] ;
wire \u_lsu.pmem[4779] ;
wire \u_lsu.pmem[4780] ;
wire \u_lsu.pmem[4781] ;
wire \u_lsu.pmem[4782] ;
wire \u_lsu.pmem[4783] ;
wire \u_lsu.pmem[4784] ;
wire \u_lsu.pmem[4785] ;
wire \u_lsu.pmem[4786] ;
wire \u_lsu.pmem[4787] ;
wire \u_lsu.pmem[4788] ;
wire \u_lsu.pmem[4789] ;
wire \u_lsu.pmem[4790] ;
wire \u_lsu.pmem[4791] ;
wire \u_lsu.pmem[4792] ;
wire \u_lsu.pmem[4793] ;
wire \u_lsu.pmem[4794] ;
wire \u_lsu.pmem[4795] ;
wire \u_lsu.pmem[4796] ;
wire \u_lsu.pmem[4797] ;
wire \u_lsu.pmem[4798] ;
wire \u_lsu.pmem[4799] ;
wire \u_lsu.pmem[4800] ;
wire \u_lsu.pmem[4801] ;
wire \u_lsu.pmem[4802] ;
wire \u_lsu.pmem[4803] ;
wire \u_lsu.pmem[4804] ;
wire \u_lsu.pmem[4805] ;
wire \u_lsu.pmem[4806] ;
wire \u_lsu.pmem[4807] ;
wire \u_lsu.pmem[4808] ;
wire \u_lsu.pmem[4809] ;
wire \u_lsu.pmem[4810] ;
wire \u_lsu.pmem[4811] ;
wire \u_lsu.pmem[4812] ;
wire \u_lsu.pmem[4813] ;
wire \u_lsu.pmem[4814] ;
wire \u_lsu.pmem[4815] ;
wire \u_lsu.pmem[4816] ;
wire \u_lsu.pmem[4817] ;
wire \u_lsu.pmem[4818] ;
wire \u_lsu.pmem[4819] ;
wire \u_lsu.pmem[4820] ;
wire \u_lsu.pmem[4821] ;
wire \u_lsu.pmem[4822] ;
wire \u_lsu.pmem[4823] ;
wire \u_lsu.pmem[4824] ;
wire \u_lsu.pmem[4825] ;
wire \u_lsu.pmem[4826] ;
wire \u_lsu.pmem[4827] ;
wire \u_lsu.pmem[4828] ;
wire \u_lsu.pmem[4829] ;
wire \u_lsu.pmem[4830] ;
wire \u_lsu.pmem[4831] ;
wire \u_lsu.pmem[4832] ;
wire \u_lsu.pmem[4833] ;
wire \u_lsu.pmem[4834] ;
wire \u_lsu.pmem[4835] ;
wire \u_lsu.pmem[4836] ;
wire \u_lsu.pmem[4837] ;
wire \u_lsu.pmem[4838] ;
wire \u_lsu.pmem[4839] ;
wire \u_lsu.pmem[4840] ;
wire \u_lsu.pmem[4841] ;
wire \u_lsu.pmem[4842] ;
wire \u_lsu.pmem[4843] ;
wire \u_lsu.pmem[4844] ;
wire \u_lsu.pmem[4845] ;
wire \u_lsu.pmem[4846] ;
wire \u_lsu.pmem[4847] ;
wire \u_lsu.pmem[4848] ;
wire \u_lsu.pmem[4849] ;
wire \u_lsu.pmem[4850] ;
wire \u_lsu.pmem[4851] ;
wire \u_lsu.pmem[4852] ;
wire \u_lsu.pmem[4853] ;
wire \u_lsu.pmem[4854] ;
wire \u_lsu.pmem[4855] ;
wire \u_lsu.pmem[4856] ;
wire \u_lsu.pmem[4857] ;
wire \u_lsu.pmem[4858] ;
wire \u_lsu.pmem[4859] ;
wire \u_lsu.pmem[4860] ;
wire \u_lsu.pmem[4861] ;
wire \u_lsu.pmem[4862] ;
wire \u_lsu.pmem[4863] ;
wire \u_lsu.pmem[4864] ;
wire \u_lsu.pmem[4865] ;
wire \u_lsu.pmem[4866] ;
wire \u_lsu.pmem[4867] ;
wire \u_lsu.pmem[4868] ;
wire \u_lsu.pmem[4869] ;
wire \u_lsu.pmem[4870] ;
wire \u_lsu.pmem[4871] ;
wire \u_lsu.pmem[4872] ;
wire \u_lsu.pmem[4873] ;
wire \u_lsu.pmem[4874] ;
wire \u_lsu.pmem[4875] ;
wire \u_lsu.pmem[4876] ;
wire \u_lsu.pmem[4877] ;
wire \u_lsu.pmem[4878] ;
wire \u_lsu.pmem[4879] ;
wire \u_lsu.pmem[4880] ;
wire \u_lsu.pmem[4881] ;
wire \u_lsu.pmem[4882] ;
wire \u_lsu.pmem[4883] ;
wire \u_lsu.pmem[4884] ;
wire \u_lsu.pmem[4885] ;
wire \u_lsu.pmem[4886] ;
wire \u_lsu.pmem[4887] ;
wire \u_lsu.pmem[4888] ;
wire \u_lsu.pmem[4889] ;
wire \u_lsu.pmem[4890] ;
wire \u_lsu.pmem[4891] ;
wire \u_lsu.pmem[4892] ;
wire \u_lsu.pmem[4893] ;
wire \u_lsu.pmem[4894] ;
wire \u_lsu.pmem[4895] ;
wire \u_lsu.pmem[4896] ;
wire \u_lsu.pmem[4897] ;
wire \u_lsu.pmem[4898] ;
wire \u_lsu.pmem[4899] ;
wire \u_lsu.pmem[4900] ;
wire \u_lsu.pmem[4901] ;
wire \u_lsu.pmem[4902] ;
wire \u_lsu.pmem[4903] ;
wire \u_lsu.pmem[4904] ;
wire \u_lsu.pmem[4905] ;
wire \u_lsu.pmem[4906] ;
wire \u_lsu.pmem[4907] ;
wire \u_lsu.pmem[4908] ;
wire \u_lsu.pmem[4909] ;
wire \u_lsu.pmem[4910] ;
wire \u_lsu.pmem[4911] ;
wire \u_lsu.pmem[4912] ;
wire \u_lsu.pmem[4913] ;
wire \u_lsu.pmem[4914] ;
wire \u_lsu.pmem[4915] ;
wire \u_lsu.pmem[4916] ;
wire \u_lsu.pmem[4917] ;
wire \u_lsu.pmem[4918] ;
wire \u_lsu.pmem[4919] ;
wire \u_lsu.pmem[4920] ;
wire \u_lsu.pmem[4921] ;
wire \u_lsu.pmem[4922] ;
wire \u_lsu.pmem[4923] ;
wire \u_lsu.pmem[4924] ;
wire \u_lsu.pmem[4925] ;
wire \u_lsu.pmem[4926] ;
wire \u_lsu.pmem[4927] ;
wire \u_lsu.pmem[4928] ;
wire \u_lsu.pmem[4929] ;
wire \u_lsu.pmem[4930] ;
wire \u_lsu.pmem[4931] ;
wire \u_lsu.pmem[4932] ;
wire \u_lsu.pmem[4933] ;
wire \u_lsu.pmem[4934] ;
wire \u_lsu.pmem[4935] ;
wire \u_lsu.pmem[4936] ;
wire \u_lsu.pmem[4937] ;
wire \u_lsu.pmem[4938] ;
wire \u_lsu.pmem[4939] ;
wire \u_lsu.pmem[4940] ;
wire \u_lsu.pmem[4941] ;
wire \u_lsu.pmem[4942] ;
wire \u_lsu.pmem[4943] ;
wire \u_lsu.pmem[4944] ;
wire \u_lsu.pmem[4945] ;
wire \u_lsu.pmem[4946] ;
wire \u_lsu.pmem[4947] ;
wire \u_lsu.pmem[4948] ;
wire \u_lsu.pmem[4949] ;
wire \u_lsu.pmem[4950] ;
wire \u_lsu.pmem[4951] ;
wire \u_lsu.pmem[4952] ;
wire \u_lsu.pmem[4953] ;
wire \u_lsu.pmem[4954] ;
wire \u_lsu.pmem[4955] ;
wire \u_lsu.pmem[4956] ;
wire \u_lsu.pmem[4957] ;
wire \u_lsu.pmem[4958] ;
wire \u_lsu.pmem[4959] ;
wire \u_lsu.pmem[4960] ;
wire \u_lsu.pmem[4961] ;
wire \u_lsu.pmem[4962] ;
wire \u_lsu.pmem[4963] ;
wire \u_lsu.pmem[4964] ;
wire \u_lsu.pmem[4965] ;
wire \u_lsu.pmem[4966] ;
wire \u_lsu.pmem[4967] ;
wire \u_lsu.pmem[4968] ;
wire \u_lsu.pmem[4969] ;
wire \u_lsu.pmem[4970] ;
wire \u_lsu.pmem[4971] ;
wire \u_lsu.pmem[4972] ;
wire \u_lsu.pmem[4973] ;
wire \u_lsu.pmem[4974] ;
wire \u_lsu.pmem[4975] ;
wire \u_lsu.pmem[4976] ;
wire \u_lsu.pmem[4977] ;
wire \u_lsu.pmem[4978] ;
wire \u_lsu.pmem[4979] ;
wire \u_lsu.pmem[4980] ;
wire \u_lsu.pmem[4981] ;
wire \u_lsu.pmem[4982] ;
wire \u_lsu.pmem[4983] ;
wire \u_lsu.pmem[4984] ;
wire \u_lsu.pmem[4985] ;
wire \u_lsu.pmem[4986] ;
wire \u_lsu.pmem[4987] ;
wire \u_lsu.pmem[4988] ;
wire \u_lsu.pmem[4989] ;
wire \u_lsu.pmem[4990] ;
wire \u_lsu.pmem[4991] ;
wire \u_lsu.pmem[4992] ;
wire \u_lsu.pmem[4993] ;
wire \u_lsu.pmem[4994] ;
wire \u_lsu.pmem[4995] ;
wire \u_lsu.pmem[4996] ;
wire \u_lsu.pmem[4997] ;
wire \u_lsu.pmem[4998] ;
wire \u_lsu.pmem[4999] ;
wire \u_lsu.pmem[5000] ;
wire \u_lsu.pmem[5001] ;
wire \u_lsu.pmem[5002] ;
wire \u_lsu.pmem[5003] ;
wire \u_lsu.pmem[5004] ;
wire \u_lsu.pmem[5005] ;
wire \u_lsu.pmem[5006] ;
wire \u_lsu.pmem[5007] ;
wire \u_lsu.pmem[5008] ;
wire \u_lsu.pmem[5009] ;
wire \u_lsu.pmem[5010] ;
wire \u_lsu.pmem[5011] ;
wire \u_lsu.pmem[5012] ;
wire \u_lsu.pmem[5013] ;
wire \u_lsu.pmem[5014] ;
wire \u_lsu.pmem[5015] ;
wire \u_lsu.pmem[5016] ;
wire \u_lsu.pmem[5017] ;
wire \u_lsu.pmem[5018] ;
wire \u_lsu.pmem[5019] ;
wire \u_lsu.pmem[5020] ;
wire \u_lsu.pmem[5021] ;
wire \u_lsu.pmem[5022] ;
wire \u_lsu.pmem[5023] ;
wire \u_lsu.pmem[5024] ;
wire \u_lsu.pmem[5025] ;
wire \u_lsu.pmem[5026] ;
wire \u_lsu.pmem[5027] ;
wire \u_lsu.pmem[5028] ;
wire \u_lsu.pmem[5029] ;
wire \u_lsu.pmem[5030] ;
wire \u_lsu.pmem[5031] ;
wire \u_lsu.pmem[5032] ;
wire \u_lsu.pmem[5033] ;
wire \u_lsu.pmem[5034] ;
wire \u_lsu.pmem[5035] ;
wire \u_lsu.pmem[5036] ;
wire \u_lsu.pmem[5037] ;
wire \u_lsu.pmem[5038] ;
wire \u_lsu.pmem[5039] ;
wire \u_lsu.pmem[5040] ;
wire \u_lsu.pmem[5041] ;
wire \u_lsu.pmem[5042] ;
wire \u_lsu.pmem[5043] ;
wire \u_lsu.pmem[5044] ;
wire \u_lsu.pmem[5045] ;
wire \u_lsu.pmem[5046] ;
wire \u_lsu.pmem[5047] ;
wire \u_lsu.pmem[5048] ;
wire \u_lsu.pmem[5049] ;
wire \u_lsu.pmem[5050] ;
wire \u_lsu.pmem[5051] ;
wire \u_lsu.pmem[5052] ;
wire \u_lsu.pmem[5053] ;
wire \u_lsu.pmem[5054] ;
wire \u_lsu.pmem[5055] ;
wire \u_lsu.pmem[5056] ;
wire \u_lsu.pmem[5057] ;
wire \u_lsu.pmem[5058] ;
wire \u_lsu.pmem[5059] ;
wire \u_lsu.pmem[5060] ;
wire \u_lsu.pmem[5061] ;
wire \u_lsu.pmem[5062] ;
wire \u_lsu.pmem[5063] ;
wire \u_lsu.pmem[5064] ;
wire \u_lsu.pmem[5065] ;
wire \u_lsu.pmem[5066] ;
wire \u_lsu.pmem[5067] ;
wire \u_lsu.pmem[5068] ;
wire \u_lsu.pmem[5069] ;
wire \u_lsu.pmem[5070] ;
wire \u_lsu.pmem[5071] ;
wire \u_lsu.pmem[5072] ;
wire \u_lsu.pmem[5073] ;
wire \u_lsu.pmem[5074] ;
wire \u_lsu.pmem[5075] ;
wire \u_lsu.pmem[5076] ;
wire \u_lsu.pmem[5077] ;
wire \u_lsu.pmem[5078] ;
wire \u_lsu.pmem[5079] ;
wire \u_lsu.pmem[5080] ;
wire \u_lsu.pmem[5081] ;
wire \u_lsu.pmem[5082] ;
wire \u_lsu.pmem[5083] ;
wire \u_lsu.pmem[5084] ;
wire \u_lsu.pmem[5085] ;
wire \u_lsu.pmem[5086] ;
wire \u_lsu.pmem[5087] ;
wire \u_lsu.pmem[5088] ;
wire \u_lsu.pmem[5089] ;
wire \u_lsu.pmem[5090] ;
wire \u_lsu.pmem[5091] ;
wire \u_lsu.pmem[5092] ;
wire \u_lsu.pmem[5093] ;
wire \u_lsu.pmem[5094] ;
wire \u_lsu.pmem[5095] ;
wire \u_lsu.pmem[5096] ;
wire \u_lsu.pmem[5097] ;
wire \u_lsu.pmem[5098] ;
wire \u_lsu.pmem[5099] ;
wire \u_lsu.pmem[5100] ;
wire \u_lsu.pmem[5101] ;
wire \u_lsu.pmem[5102] ;
wire \u_lsu.pmem[5103] ;
wire \u_lsu.pmem[5104] ;
wire \u_lsu.pmem[5105] ;
wire \u_lsu.pmem[5106] ;
wire \u_lsu.pmem[5107] ;
wire \u_lsu.pmem[5108] ;
wire \u_lsu.pmem[5109] ;
wire \u_lsu.pmem[5110] ;
wire \u_lsu.pmem[5111] ;
wire \u_lsu.pmem[5112] ;
wire \u_lsu.pmem[5113] ;
wire \u_lsu.pmem[5114] ;
wire \u_lsu.pmem[5115] ;
wire \u_lsu.pmem[5116] ;
wire \u_lsu.pmem[5117] ;
wire \u_lsu.pmem[5118] ;
wire \u_lsu.pmem[5119] ;
wire \u_lsu.pmem[5120] ;
wire \u_lsu.pmem[5121] ;
wire \u_lsu.pmem[5122] ;
wire \u_lsu.pmem[5123] ;
wire \u_lsu.pmem[5124] ;
wire \u_lsu.pmem[5125] ;
wire \u_lsu.pmem[5126] ;
wire \u_lsu.pmem[5127] ;
wire \u_lsu.pmem[5128] ;
wire \u_lsu.pmem[5129] ;
wire \u_lsu.pmem[5130] ;
wire \u_lsu.pmem[5131] ;
wire \u_lsu.pmem[5132] ;
wire \u_lsu.pmem[5133] ;
wire \u_lsu.pmem[5134] ;
wire \u_lsu.pmem[5135] ;
wire \u_lsu.pmem[5136] ;
wire \u_lsu.pmem[5137] ;
wire \u_lsu.pmem[5138] ;
wire \u_lsu.pmem[5139] ;
wire \u_lsu.pmem[5140] ;
wire \u_lsu.pmem[5141] ;
wire \u_lsu.pmem[5142] ;
wire \u_lsu.pmem[5143] ;
wire \u_lsu.pmem[5144] ;
wire \u_lsu.pmem[5145] ;
wire \u_lsu.pmem[5146] ;
wire \u_lsu.pmem[5147] ;
wire \u_lsu.pmem[5148] ;
wire \u_lsu.pmem[5149] ;
wire \u_lsu.pmem[5150] ;
wire \u_lsu.pmem[5151] ;
wire \u_lsu.pmem[5152] ;
wire \u_lsu.pmem[5153] ;
wire \u_lsu.pmem[5154] ;
wire \u_lsu.pmem[5155] ;
wire \u_lsu.pmem[5156] ;
wire \u_lsu.pmem[5157] ;
wire \u_lsu.pmem[5158] ;
wire \u_lsu.pmem[5159] ;
wire \u_lsu.pmem[5160] ;
wire \u_lsu.pmem[5161] ;
wire \u_lsu.pmem[5162] ;
wire \u_lsu.pmem[5163] ;
wire \u_lsu.pmem[5164] ;
wire \u_lsu.pmem[5165] ;
wire \u_lsu.pmem[5166] ;
wire \u_lsu.pmem[5167] ;
wire \u_lsu.pmem[5168] ;
wire \u_lsu.pmem[5169] ;
wire \u_lsu.pmem[5170] ;
wire \u_lsu.pmem[5171] ;
wire \u_lsu.pmem[5172] ;
wire \u_lsu.pmem[5173] ;
wire \u_lsu.pmem[5174] ;
wire \u_lsu.pmem[5175] ;
wire \u_lsu.pmem[5176] ;
wire \u_lsu.pmem[5177] ;
wire \u_lsu.pmem[5178] ;
wire \u_lsu.pmem[5179] ;
wire \u_lsu.pmem[5180] ;
wire \u_lsu.pmem[5181] ;
wire \u_lsu.pmem[5182] ;
wire \u_lsu.pmem[5183] ;
wire \u_lsu.pmem[5184] ;
wire \u_lsu.pmem[5185] ;
wire \u_lsu.pmem[5186] ;
wire \u_lsu.pmem[5187] ;
wire \u_lsu.pmem[5188] ;
wire \u_lsu.pmem[5189] ;
wire \u_lsu.pmem[5190] ;
wire \u_lsu.pmem[5191] ;
wire \u_lsu.pmem[5192] ;
wire \u_lsu.pmem[5193] ;
wire \u_lsu.pmem[5194] ;
wire \u_lsu.pmem[5195] ;
wire \u_lsu.pmem[5196] ;
wire \u_lsu.pmem[5197] ;
wire \u_lsu.pmem[5198] ;
wire \u_lsu.pmem[5199] ;
wire \u_lsu.pmem[5200] ;
wire \u_lsu.pmem[5201] ;
wire \u_lsu.pmem[5202] ;
wire \u_lsu.pmem[5203] ;
wire \u_lsu.pmem[5204] ;
wire \u_lsu.pmem[5205] ;
wire \u_lsu.pmem[5206] ;
wire \u_lsu.pmem[5207] ;
wire \u_lsu.pmem[5208] ;
wire \u_lsu.pmem[5209] ;
wire \u_lsu.pmem[5210] ;
wire \u_lsu.pmem[5211] ;
wire \u_lsu.pmem[5212] ;
wire \u_lsu.pmem[5213] ;
wire \u_lsu.pmem[5214] ;
wire \u_lsu.pmem[5215] ;
wire \u_lsu.pmem[5216] ;
wire \u_lsu.pmem[5217] ;
wire \u_lsu.pmem[5218] ;
wire \u_lsu.pmem[5219] ;
wire \u_lsu.pmem[5220] ;
wire \u_lsu.pmem[5221] ;
wire \u_lsu.pmem[5222] ;
wire \u_lsu.pmem[5223] ;
wire \u_lsu.pmem[5224] ;
wire \u_lsu.pmem[5225] ;
wire \u_lsu.pmem[5226] ;
wire \u_lsu.pmem[5227] ;
wire \u_lsu.pmem[5228] ;
wire \u_lsu.pmem[5229] ;
wire \u_lsu.pmem[5230] ;
wire \u_lsu.pmem[5231] ;
wire \u_lsu.pmem[5232] ;
wire \u_lsu.pmem[5233] ;
wire \u_lsu.pmem[5234] ;
wire \u_lsu.pmem[5235] ;
wire \u_lsu.pmem[5236] ;
wire \u_lsu.pmem[5237] ;
wire \u_lsu.pmem[5238] ;
wire \u_lsu.pmem[5239] ;
wire \u_lsu.pmem[5240] ;
wire \u_lsu.pmem[5241] ;
wire \u_lsu.pmem[5242] ;
wire \u_lsu.pmem[5243] ;
wire \u_lsu.pmem[5244] ;
wire \u_lsu.pmem[5245] ;
wire \u_lsu.pmem[5246] ;
wire \u_lsu.pmem[5247] ;
wire \u_lsu.pmem[5248] ;
wire \u_lsu.pmem[5249] ;
wire \u_lsu.pmem[5250] ;
wire \u_lsu.pmem[5251] ;
wire \u_lsu.pmem[5252] ;
wire \u_lsu.pmem[5253] ;
wire \u_lsu.pmem[5254] ;
wire \u_lsu.pmem[5255] ;
wire \u_lsu.pmem[5256] ;
wire \u_lsu.pmem[5257] ;
wire \u_lsu.pmem[5258] ;
wire \u_lsu.pmem[5259] ;
wire \u_lsu.pmem[5260] ;
wire \u_lsu.pmem[5261] ;
wire \u_lsu.pmem[5262] ;
wire \u_lsu.pmem[5263] ;
wire \u_lsu.pmem[5264] ;
wire \u_lsu.pmem[5265] ;
wire \u_lsu.pmem[5266] ;
wire \u_lsu.pmem[5267] ;
wire \u_lsu.pmem[5268] ;
wire \u_lsu.pmem[5269] ;
wire \u_lsu.pmem[5270] ;
wire \u_lsu.pmem[5271] ;
wire \u_lsu.pmem[5272] ;
wire \u_lsu.pmem[5273] ;
wire \u_lsu.pmem[5274] ;
wire \u_lsu.pmem[5275] ;
wire \u_lsu.pmem[5276] ;
wire \u_lsu.pmem[5277] ;
wire \u_lsu.pmem[5278] ;
wire \u_lsu.pmem[5279] ;
wire \u_lsu.pmem[5280] ;
wire \u_lsu.pmem[5281] ;
wire \u_lsu.pmem[5282] ;
wire \u_lsu.pmem[5283] ;
wire \u_lsu.pmem[5284] ;
wire \u_lsu.pmem[5285] ;
wire \u_lsu.pmem[5286] ;
wire \u_lsu.pmem[5287] ;
wire \u_lsu.pmem[5288] ;
wire \u_lsu.pmem[5289] ;
wire \u_lsu.pmem[5290] ;
wire \u_lsu.pmem[5291] ;
wire \u_lsu.pmem[5292] ;
wire \u_lsu.pmem[5293] ;
wire \u_lsu.pmem[5294] ;
wire \u_lsu.pmem[5295] ;
wire \u_lsu.pmem[5296] ;
wire \u_lsu.pmem[5297] ;
wire \u_lsu.pmem[5298] ;
wire \u_lsu.pmem[5299] ;
wire \u_lsu.pmem[5300] ;
wire \u_lsu.pmem[5301] ;
wire \u_lsu.pmem[5302] ;
wire \u_lsu.pmem[5303] ;
wire \u_lsu.pmem[5304] ;
wire \u_lsu.pmem[5305] ;
wire \u_lsu.pmem[5306] ;
wire \u_lsu.pmem[5307] ;
wire \u_lsu.pmem[5308] ;
wire \u_lsu.pmem[5309] ;
wire \u_lsu.pmem[5310] ;
wire \u_lsu.pmem[5311] ;
wire \u_lsu.pmem[5312] ;
wire \u_lsu.pmem[5313] ;
wire \u_lsu.pmem[5314] ;
wire \u_lsu.pmem[5315] ;
wire \u_lsu.pmem[5316] ;
wire \u_lsu.pmem[5317] ;
wire \u_lsu.pmem[5318] ;
wire \u_lsu.pmem[5319] ;
wire \u_lsu.pmem[5320] ;
wire \u_lsu.pmem[5321] ;
wire \u_lsu.pmem[5322] ;
wire \u_lsu.pmem[5323] ;
wire \u_lsu.pmem[5324] ;
wire \u_lsu.pmem[5325] ;
wire \u_lsu.pmem[5326] ;
wire \u_lsu.pmem[5327] ;
wire \u_lsu.pmem[5328] ;
wire \u_lsu.pmem[5329] ;
wire \u_lsu.pmem[5330] ;
wire \u_lsu.pmem[5331] ;
wire \u_lsu.pmem[5332] ;
wire \u_lsu.pmem[5333] ;
wire \u_lsu.pmem[5334] ;
wire \u_lsu.pmem[5335] ;
wire \u_lsu.pmem[5336] ;
wire \u_lsu.pmem[5337] ;
wire \u_lsu.pmem[5338] ;
wire \u_lsu.pmem[5339] ;
wire \u_lsu.pmem[5340] ;
wire \u_lsu.pmem[5341] ;
wire \u_lsu.pmem[5342] ;
wire \u_lsu.pmem[5343] ;
wire \u_lsu.pmem[5344] ;
wire \u_lsu.pmem[5345] ;
wire \u_lsu.pmem[5346] ;
wire \u_lsu.pmem[5347] ;
wire \u_lsu.pmem[5348] ;
wire \u_lsu.pmem[5349] ;
wire \u_lsu.pmem[5350] ;
wire \u_lsu.pmem[5351] ;
wire \u_lsu.pmem[5352] ;
wire \u_lsu.pmem[5353] ;
wire \u_lsu.pmem[5354] ;
wire \u_lsu.pmem[5355] ;
wire \u_lsu.pmem[5356] ;
wire \u_lsu.pmem[5357] ;
wire \u_lsu.pmem[5358] ;
wire \u_lsu.pmem[5359] ;
wire \u_lsu.pmem[5360] ;
wire \u_lsu.pmem[5361] ;
wire \u_lsu.pmem[5362] ;
wire \u_lsu.pmem[5363] ;
wire \u_lsu.pmem[5364] ;
wire \u_lsu.pmem[5365] ;
wire \u_lsu.pmem[5366] ;
wire \u_lsu.pmem[5367] ;
wire \u_lsu.pmem[5368] ;
wire \u_lsu.pmem[5369] ;
wire \u_lsu.pmem[5370] ;
wire \u_lsu.pmem[5371] ;
wire \u_lsu.pmem[5372] ;
wire \u_lsu.pmem[5373] ;
wire \u_lsu.pmem[5374] ;
wire \u_lsu.pmem[5375] ;
wire \u_lsu.pmem[5376] ;
wire \u_lsu.pmem[5377] ;
wire \u_lsu.pmem[5378] ;
wire \u_lsu.pmem[5379] ;
wire \u_lsu.pmem[5380] ;
wire \u_lsu.pmem[5381] ;
wire \u_lsu.pmem[5382] ;
wire \u_lsu.pmem[5383] ;
wire \u_lsu.pmem[5384] ;
wire \u_lsu.pmem[5385] ;
wire \u_lsu.pmem[5386] ;
wire \u_lsu.pmem[5387] ;
wire \u_lsu.pmem[5388] ;
wire \u_lsu.pmem[5389] ;
wire \u_lsu.pmem[5390] ;
wire \u_lsu.pmem[5391] ;
wire \u_lsu.pmem[5392] ;
wire \u_lsu.pmem[5393] ;
wire \u_lsu.pmem[5394] ;
wire \u_lsu.pmem[5395] ;
wire \u_lsu.pmem[5396] ;
wire \u_lsu.pmem[5397] ;
wire \u_lsu.pmem[5398] ;
wire \u_lsu.pmem[5399] ;
wire \u_lsu.pmem[5400] ;
wire \u_lsu.pmem[5401] ;
wire \u_lsu.pmem[5402] ;
wire \u_lsu.pmem[5403] ;
wire \u_lsu.pmem[5404] ;
wire \u_lsu.pmem[5405] ;
wire \u_lsu.pmem[5406] ;
wire \u_lsu.pmem[5407] ;
wire \u_lsu.pmem[5408] ;
wire \u_lsu.pmem[5409] ;
wire \u_lsu.pmem[5410] ;
wire \u_lsu.pmem[5411] ;
wire \u_lsu.pmem[5412] ;
wire \u_lsu.pmem[5413] ;
wire \u_lsu.pmem[5414] ;
wire \u_lsu.pmem[5415] ;
wire \u_lsu.pmem[5416] ;
wire \u_lsu.pmem[5417] ;
wire \u_lsu.pmem[5418] ;
wire \u_lsu.pmem[5419] ;
wire \u_lsu.pmem[5420] ;
wire \u_lsu.pmem[5421] ;
wire \u_lsu.pmem[5422] ;
wire \u_lsu.pmem[5423] ;
wire \u_lsu.pmem[5424] ;
wire \u_lsu.pmem[5425] ;
wire \u_lsu.pmem[5426] ;
wire \u_lsu.pmem[5427] ;
wire \u_lsu.pmem[5428] ;
wire \u_lsu.pmem[5429] ;
wire \u_lsu.pmem[5430] ;
wire \u_lsu.pmem[5431] ;
wire \u_lsu.pmem[5432] ;
wire \u_lsu.pmem[5433] ;
wire \u_lsu.pmem[5434] ;
wire \u_lsu.pmem[5435] ;
wire \u_lsu.pmem[5436] ;
wire \u_lsu.pmem[5437] ;
wire \u_lsu.pmem[5438] ;
wire \u_lsu.pmem[5439] ;
wire \u_lsu.pmem[5440] ;
wire \u_lsu.pmem[5441] ;
wire \u_lsu.pmem[5442] ;
wire \u_lsu.pmem[5443] ;
wire \u_lsu.pmem[5444] ;
wire \u_lsu.pmem[5445] ;
wire \u_lsu.pmem[5446] ;
wire \u_lsu.pmem[5447] ;
wire \u_lsu.pmem[5448] ;
wire \u_lsu.pmem[5449] ;
wire \u_lsu.pmem[5450] ;
wire \u_lsu.pmem[5451] ;
wire \u_lsu.pmem[5452] ;
wire \u_lsu.pmem[5453] ;
wire \u_lsu.pmem[5454] ;
wire \u_lsu.pmem[5455] ;
wire \u_lsu.pmem[5456] ;
wire \u_lsu.pmem[5457] ;
wire \u_lsu.pmem[5458] ;
wire \u_lsu.pmem[5459] ;
wire \u_lsu.pmem[5460] ;
wire \u_lsu.pmem[5461] ;
wire \u_lsu.pmem[5462] ;
wire \u_lsu.pmem[5463] ;
wire \u_lsu.pmem[5464] ;
wire \u_lsu.pmem[5465] ;
wire \u_lsu.pmem[5466] ;
wire \u_lsu.pmem[5467] ;
wire \u_lsu.pmem[5468] ;
wire \u_lsu.pmem[5469] ;
wire \u_lsu.pmem[5470] ;
wire \u_lsu.pmem[5471] ;
wire \u_lsu.pmem[5472] ;
wire \u_lsu.pmem[5473] ;
wire \u_lsu.pmem[5474] ;
wire \u_lsu.pmem[5475] ;
wire \u_lsu.pmem[5476] ;
wire \u_lsu.pmem[5477] ;
wire \u_lsu.pmem[5478] ;
wire \u_lsu.pmem[5479] ;
wire \u_lsu.pmem[5480] ;
wire \u_lsu.pmem[5481] ;
wire \u_lsu.pmem[5482] ;
wire \u_lsu.pmem[5483] ;
wire \u_lsu.pmem[5484] ;
wire \u_lsu.pmem[5485] ;
wire \u_lsu.pmem[5486] ;
wire \u_lsu.pmem[5487] ;
wire \u_lsu.pmem[5488] ;
wire \u_lsu.pmem[5489] ;
wire \u_lsu.pmem[5490] ;
wire \u_lsu.pmem[5491] ;
wire \u_lsu.pmem[5492] ;
wire \u_lsu.pmem[5493] ;
wire \u_lsu.pmem[5494] ;
wire \u_lsu.pmem[5495] ;
wire \u_lsu.pmem[5496] ;
wire \u_lsu.pmem[5497] ;
wire \u_lsu.pmem[5498] ;
wire \u_lsu.pmem[5499] ;
wire \u_lsu.pmem[5500] ;
wire \u_lsu.pmem[5501] ;
wire \u_lsu.pmem[5502] ;
wire \u_lsu.pmem[5503] ;
wire \u_lsu.pmem[5504] ;
wire \u_lsu.pmem[5505] ;
wire \u_lsu.pmem[5506] ;
wire \u_lsu.pmem[5507] ;
wire \u_lsu.pmem[5508] ;
wire \u_lsu.pmem[5509] ;
wire \u_lsu.pmem[5510] ;
wire \u_lsu.pmem[5511] ;
wire \u_lsu.pmem[5512] ;
wire \u_lsu.pmem[5513] ;
wire \u_lsu.pmem[5514] ;
wire \u_lsu.pmem[5515] ;
wire \u_lsu.pmem[5516] ;
wire \u_lsu.pmem[5517] ;
wire \u_lsu.pmem[5518] ;
wire \u_lsu.pmem[5519] ;
wire \u_lsu.pmem[5520] ;
wire \u_lsu.pmem[5521] ;
wire \u_lsu.pmem[5522] ;
wire \u_lsu.pmem[5523] ;
wire \u_lsu.pmem[5524] ;
wire \u_lsu.pmem[5525] ;
wire \u_lsu.pmem[5526] ;
wire \u_lsu.pmem[5527] ;
wire \u_lsu.pmem[5528] ;
wire \u_lsu.pmem[5529] ;
wire \u_lsu.pmem[5530] ;
wire \u_lsu.pmem[5531] ;
wire \u_lsu.pmem[5532] ;
wire \u_lsu.pmem[5533] ;
wire \u_lsu.pmem[5534] ;
wire \u_lsu.pmem[5535] ;
wire \u_lsu.pmem[5536] ;
wire \u_lsu.pmem[5537] ;
wire \u_lsu.pmem[5538] ;
wire \u_lsu.pmem[5539] ;
wire \u_lsu.pmem[5540] ;
wire \u_lsu.pmem[5541] ;
wire \u_lsu.pmem[5542] ;
wire \u_lsu.pmem[5543] ;
wire \u_lsu.pmem[5544] ;
wire \u_lsu.pmem[5545] ;
wire \u_lsu.pmem[5546] ;
wire \u_lsu.pmem[5547] ;
wire \u_lsu.pmem[5548] ;
wire \u_lsu.pmem[5549] ;
wire \u_lsu.pmem[5550] ;
wire \u_lsu.pmem[5551] ;
wire \u_lsu.pmem[5552] ;
wire \u_lsu.pmem[5553] ;
wire \u_lsu.pmem[5554] ;
wire \u_lsu.pmem[5555] ;
wire \u_lsu.pmem[5556] ;
wire \u_lsu.pmem[5557] ;
wire \u_lsu.pmem[5558] ;
wire \u_lsu.pmem[5559] ;
wire \u_lsu.pmem[5560] ;
wire \u_lsu.pmem[5561] ;
wire \u_lsu.pmem[5562] ;
wire \u_lsu.pmem[5563] ;
wire \u_lsu.pmem[5564] ;
wire \u_lsu.pmem[5565] ;
wire \u_lsu.pmem[5566] ;
wire \u_lsu.pmem[5567] ;
wire \u_lsu.pmem[5568] ;
wire \u_lsu.pmem[5569] ;
wire \u_lsu.pmem[5570] ;
wire \u_lsu.pmem[5571] ;
wire \u_lsu.pmem[5572] ;
wire \u_lsu.pmem[5573] ;
wire \u_lsu.pmem[5574] ;
wire \u_lsu.pmem[5575] ;
wire \u_lsu.pmem[5576] ;
wire \u_lsu.pmem[5577] ;
wire \u_lsu.pmem[5578] ;
wire \u_lsu.pmem[5579] ;
wire \u_lsu.pmem[5580] ;
wire \u_lsu.pmem[5581] ;
wire \u_lsu.pmem[5582] ;
wire \u_lsu.pmem[5583] ;
wire \u_lsu.pmem[5584] ;
wire \u_lsu.pmem[5585] ;
wire \u_lsu.pmem[5586] ;
wire \u_lsu.pmem[5587] ;
wire \u_lsu.pmem[5588] ;
wire \u_lsu.pmem[5589] ;
wire \u_lsu.pmem[5590] ;
wire \u_lsu.pmem[5591] ;
wire \u_lsu.pmem[5592] ;
wire \u_lsu.pmem[5593] ;
wire \u_lsu.pmem[5594] ;
wire \u_lsu.pmem[5595] ;
wire \u_lsu.pmem[5596] ;
wire \u_lsu.pmem[5597] ;
wire \u_lsu.pmem[5598] ;
wire \u_lsu.pmem[5599] ;
wire \u_lsu.pmem[5600] ;
wire \u_lsu.pmem[5601] ;
wire \u_lsu.pmem[5602] ;
wire \u_lsu.pmem[5603] ;
wire \u_lsu.pmem[5604] ;
wire \u_lsu.pmem[5605] ;
wire \u_lsu.pmem[5606] ;
wire \u_lsu.pmem[5607] ;
wire \u_lsu.pmem[5608] ;
wire \u_lsu.pmem[5609] ;
wire \u_lsu.pmem[5610] ;
wire \u_lsu.pmem[5611] ;
wire \u_lsu.pmem[5612] ;
wire \u_lsu.pmem[5613] ;
wire \u_lsu.pmem[5614] ;
wire \u_lsu.pmem[5615] ;
wire \u_lsu.pmem[5616] ;
wire \u_lsu.pmem[5617] ;
wire \u_lsu.pmem[5618] ;
wire \u_lsu.pmem[5619] ;
wire \u_lsu.pmem[5620] ;
wire \u_lsu.pmem[5621] ;
wire \u_lsu.pmem[5622] ;
wire \u_lsu.pmem[5623] ;
wire \u_lsu.pmem[5624] ;
wire \u_lsu.pmem[5625] ;
wire \u_lsu.pmem[5626] ;
wire \u_lsu.pmem[5627] ;
wire \u_lsu.pmem[5628] ;
wire \u_lsu.pmem[5629] ;
wire \u_lsu.pmem[5630] ;
wire \u_lsu.pmem[5631] ;
wire \u_lsu.pmem[5632] ;
wire \u_lsu.pmem[5633] ;
wire \u_lsu.pmem[5634] ;
wire \u_lsu.pmem[5635] ;
wire \u_lsu.pmem[5636] ;
wire \u_lsu.pmem[5637] ;
wire \u_lsu.pmem[5638] ;
wire \u_lsu.pmem[5639] ;
wire \u_lsu.pmem[5640] ;
wire \u_lsu.pmem[5641] ;
wire \u_lsu.pmem[5642] ;
wire \u_lsu.pmem[5643] ;
wire \u_lsu.pmem[5644] ;
wire \u_lsu.pmem[5645] ;
wire \u_lsu.pmem[5646] ;
wire \u_lsu.pmem[5647] ;
wire \u_lsu.pmem[5648] ;
wire \u_lsu.pmem[5649] ;
wire \u_lsu.pmem[5650] ;
wire \u_lsu.pmem[5651] ;
wire \u_lsu.pmem[5652] ;
wire \u_lsu.pmem[5653] ;
wire \u_lsu.pmem[5654] ;
wire \u_lsu.pmem[5655] ;
wire \u_lsu.pmem[5656] ;
wire \u_lsu.pmem[5657] ;
wire \u_lsu.pmem[5658] ;
wire \u_lsu.pmem[5659] ;
wire \u_lsu.pmem[5660] ;
wire \u_lsu.pmem[5661] ;
wire \u_lsu.pmem[5662] ;
wire \u_lsu.pmem[5663] ;
wire \u_lsu.pmem[5664] ;
wire \u_lsu.pmem[5665] ;
wire \u_lsu.pmem[5666] ;
wire \u_lsu.pmem[5667] ;
wire \u_lsu.pmem[5668] ;
wire \u_lsu.pmem[5669] ;
wire \u_lsu.pmem[5670] ;
wire \u_lsu.pmem[5671] ;
wire \u_lsu.pmem[5672] ;
wire \u_lsu.pmem[5673] ;
wire \u_lsu.pmem[5674] ;
wire \u_lsu.pmem[5675] ;
wire \u_lsu.pmem[5676] ;
wire \u_lsu.pmem[5677] ;
wire \u_lsu.pmem[5678] ;
wire \u_lsu.pmem[5679] ;
wire \u_lsu.pmem[5680] ;
wire \u_lsu.pmem[5681] ;
wire \u_lsu.pmem[5682] ;
wire \u_lsu.pmem[5683] ;
wire \u_lsu.pmem[5684] ;
wire \u_lsu.pmem[5685] ;
wire \u_lsu.pmem[5686] ;
wire \u_lsu.pmem[5687] ;
wire \u_lsu.pmem[5688] ;
wire \u_lsu.pmem[5689] ;
wire \u_lsu.pmem[5690] ;
wire \u_lsu.pmem[5691] ;
wire \u_lsu.pmem[5692] ;
wire \u_lsu.pmem[5693] ;
wire \u_lsu.pmem[5694] ;
wire \u_lsu.pmem[5695] ;
wire \u_lsu.pmem[5696] ;
wire \u_lsu.pmem[5697] ;
wire \u_lsu.pmem[5698] ;
wire \u_lsu.pmem[5699] ;
wire \u_lsu.pmem[5700] ;
wire \u_lsu.pmem[5701] ;
wire \u_lsu.pmem[5702] ;
wire \u_lsu.pmem[5703] ;
wire \u_lsu.pmem[5704] ;
wire \u_lsu.pmem[5705] ;
wire \u_lsu.pmem[5706] ;
wire \u_lsu.pmem[5707] ;
wire \u_lsu.pmem[5708] ;
wire \u_lsu.pmem[5709] ;
wire \u_lsu.pmem[5710] ;
wire \u_lsu.pmem[5711] ;
wire \u_lsu.pmem[5712] ;
wire \u_lsu.pmem[5713] ;
wire \u_lsu.pmem[5714] ;
wire \u_lsu.pmem[5715] ;
wire \u_lsu.pmem[5716] ;
wire \u_lsu.pmem[5717] ;
wire \u_lsu.pmem[5718] ;
wire \u_lsu.pmem[5719] ;
wire \u_lsu.pmem[5720] ;
wire \u_lsu.pmem[5721] ;
wire \u_lsu.pmem[5722] ;
wire \u_lsu.pmem[5723] ;
wire \u_lsu.pmem[5724] ;
wire \u_lsu.pmem[5725] ;
wire \u_lsu.pmem[5726] ;
wire \u_lsu.pmem[5727] ;
wire \u_lsu.pmem[5728] ;
wire \u_lsu.pmem[5729] ;
wire \u_lsu.pmem[5730] ;
wire \u_lsu.pmem[5731] ;
wire \u_lsu.pmem[5732] ;
wire \u_lsu.pmem[5733] ;
wire \u_lsu.pmem[5734] ;
wire \u_lsu.pmem[5735] ;
wire \u_lsu.pmem[5736] ;
wire \u_lsu.pmem[5737] ;
wire \u_lsu.pmem[5738] ;
wire \u_lsu.pmem[5739] ;
wire \u_lsu.pmem[5740] ;
wire \u_lsu.pmem[5741] ;
wire \u_lsu.pmem[5742] ;
wire \u_lsu.pmem[5743] ;
wire \u_lsu.pmem[5744] ;
wire \u_lsu.pmem[5745] ;
wire \u_lsu.pmem[5746] ;
wire \u_lsu.pmem[5747] ;
wire \u_lsu.pmem[5748] ;
wire \u_lsu.pmem[5749] ;
wire \u_lsu.pmem[5750] ;
wire \u_lsu.pmem[5751] ;
wire \u_lsu.pmem[5752] ;
wire \u_lsu.pmem[5753] ;
wire \u_lsu.pmem[5754] ;
wire \u_lsu.pmem[5755] ;
wire \u_lsu.pmem[5756] ;
wire \u_lsu.pmem[5757] ;
wire \u_lsu.pmem[5758] ;
wire \u_lsu.pmem[5759] ;
wire \u_lsu.pmem[5760] ;
wire \u_lsu.pmem[5761] ;
wire \u_lsu.pmem[5762] ;
wire \u_lsu.pmem[5763] ;
wire \u_lsu.pmem[5764] ;
wire \u_lsu.pmem[5765] ;
wire \u_lsu.pmem[5766] ;
wire \u_lsu.pmem[5767] ;
wire \u_lsu.pmem[5768] ;
wire \u_lsu.pmem[5769] ;
wire \u_lsu.pmem[5770] ;
wire \u_lsu.pmem[5771] ;
wire \u_lsu.pmem[5772] ;
wire \u_lsu.pmem[5773] ;
wire \u_lsu.pmem[5774] ;
wire \u_lsu.pmem[5775] ;
wire \u_lsu.pmem[5776] ;
wire \u_lsu.pmem[5777] ;
wire \u_lsu.pmem[5778] ;
wire \u_lsu.pmem[5779] ;
wire \u_lsu.pmem[5780] ;
wire \u_lsu.pmem[5781] ;
wire \u_lsu.pmem[5782] ;
wire \u_lsu.pmem[5783] ;
wire \u_lsu.pmem[5784] ;
wire \u_lsu.pmem[5785] ;
wire \u_lsu.pmem[5786] ;
wire \u_lsu.pmem[5787] ;
wire \u_lsu.pmem[5788] ;
wire \u_lsu.pmem[5789] ;
wire \u_lsu.pmem[5790] ;
wire \u_lsu.pmem[5791] ;
wire \u_lsu.pmem[5792] ;
wire \u_lsu.pmem[5793] ;
wire \u_lsu.pmem[5794] ;
wire \u_lsu.pmem[5795] ;
wire \u_lsu.pmem[5796] ;
wire \u_lsu.pmem[5797] ;
wire \u_lsu.pmem[5798] ;
wire \u_lsu.pmem[5799] ;
wire \u_lsu.pmem[5800] ;
wire \u_lsu.pmem[5801] ;
wire \u_lsu.pmem[5802] ;
wire \u_lsu.pmem[5803] ;
wire \u_lsu.pmem[5804] ;
wire \u_lsu.pmem[5805] ;
wire \u_lsu.pmem[5806] ;
wire \u_lsu.pmem[5807] ;
wire \u_lsu.pmem[5808] ;
wire \u_lsu.pmem[5809] ;
wire \u_lsu.pmem[5810] ;
wire \u_lsu.pmem[5811] ;
wire \u_lsu.pmem[5812] ;
wire \u_lsu.pmem[5813] ;
wire \u_lsu.pmem[5814] ;
wire \u_lsu.pmem[5815] ;
wire \u_lsu.pmem[5816] ;
wire \u_lsu.pmem[5817] ;
wire \u_lsu.pmem[5818] ;
wire \u_lsu.pmem[5819] ;
wire \u_lsu.pmem[5820] ;
wire \u_lsu.pmem[5821] ;
wire \u_lsu.pmem[5822] ;
wire \u_lsu.pmem[5823] ;
wire \u_lsu.pmem[5824] ;
wire \u_lsu.pmem[5825] ;
wire \u_lsu.pmem[5826] ;
wire \u_lsu.pmem[5827] ;
wire \u_lsu.pmem[5828] ;
wire \u_lsu.pmem[5829] ;
wire \u_lsu.pmem[5830] ;
wire \u_lsu.pmem[5831] ;
wire \u_lsu.pmem[5832] ;
wire \u_lsu.pmem[5833] ;
wire \u_lsu.pmem[5834] ;
wire \u_lsu.pmem[5835] ;
wire \u_lsu.pmem[5836] ;
wire \u_lsu.pmem[5837] ;
wire \u_lsu.pmem[5838] ;
wire \u_lsu.pmem[5839] ;
wire \u_lsu.pmem[5840] ;
wire \u_lsu.pmem[5841] ;
wire \u_lsu.pmem[5842] ;
wire \u_lsu.pmem[5843] ;
wire \u_lsu.pmem[5844] ;
wire \u_lsu.pmem[5845] ;
wire \u_lsu.pmem[5846] ;
wire \u_lsu.pmem[5847] ;
wire \u_lsu.pmem[5848] ;
wire \u_lsu.pmem[5849] ;
wire \u_lsu.pmem[5850] ;
wire \u_lsu.pmem[5851] ;
wire \u_lsu.pmem[5852] ;
wire \u_lsu.pmem[5853] ;
wire \u_lsu.pmem[5854] ;
wire \u_lsu.pmem[5855] ;
wire \u_lsu.pmem[5856] ;
wire \u_lsu.pmem[5857] ;
wire \u_lsu.pmem[5858] ;
wire \u_lsu.pmem[5859] ;
wire \u_lsu.pmem[5860] ;
wire \u_lsu.pmem[5861] ;
wire \u_lsu.pmem[5862] ;
wire \u_lsu.pmem[5863] ;
wire \u_lsu.pmem[5864] ;
wire \u_lsu.pmem[5865] ;
wire \u_lsu.pmem[5866] ;
wire \u_lsu.pmem[5867] ;
wire \u_lsu.pmem[5868] ;
wire \u_lsu.pmem[5869] ;
wire \u_lsu.pmem[5870] ;
wire \u_lsu.pmem[5871] ;
wire \u_lsu.pmem[5872] ;
wire \u_lsu.pmem[5873] ;
wire \u_lsu.pmem[5874] ;
wire \u_lsu.pmem[5875] ;
wire \u_lsu.pmem[5876] ;
wire \u_lsu.pmem[5877] ;
wire \u_lsu.pmem[5878] ;
wire \u_lsu.pmem[5879] ;
wire \u_lsu.pmem[5880] ;
wire \u_lsu.pmem[5881] ;
wire \u_lsu.pmem[5882] ;
wire \u_lsu.pmem[5883] ;
wire \u_lsu.pmem[5884] ;
wire \u_lsu.pmem[5885] ;
wire \u_lsu.pmem[5886] ;
wire \u_lsu.pmem[5887] ;
wire \u_lsu.pmem[5888] ;
wire \u_lsu.pmem[5889] ;
wire \u_lsu.pmem[5890] ;
wire \u_lsu.pmem[5891] ;
wire \u_lsu.pmem[5892] ;
wire \u_lsu.pmem[5893] ;
wire \u_lsu.pmem[5894] ;
wire \u_lsu.pmem[5895] ;
wire \u_lsu.pmem[5896] ;
wire \u_lsu.pmem[5897] ;
wire \u_lsu.pmem[5898] ;
wire \u_lsu.pmem[5899] ;
wire \u_lsu.pmem[5900] ;
wire \u_lsu.pmem[5901] ;
wire \u_lsu.pmem[5902] ;
wire \u_lsu.pmem[5903] ;
wire \u_lsu.pmem[5904] ;
wire \u_lsu.pmem[5905] ;
wire \u_lsu.pmem[5906] ;
wire \u_lsu.pmem[5907] ;
wire \u_lsu.pmem[5908] ;
wire \u_lsu.pmem[5909] ;
wire \u_lsu.pmem[5910] ;
wire \u_lsu.pmem[5911] ;
wire \u_lsu.pmem[5912] ;
wire \u_lsu.pmem[5913] ;
wire \u_lsu.pmem[5914] ;
wire \u_lsu.pmem[5915] ;
wire \u_lsu.pmem[5916] ;
wire \u_lsu.pmem[5917] ;
wire \u_lsu.pmem[5918] ;
wire \u_lsu.pmem[5919] ;
wire \u_lsu.pmem[5920] ;
wire \u_lsu.pmem[5921] ;
wire \u_lsu.pmem[5922] ;
wire \u_lsu.pmem[5923] ;
wire \u_lsu.pmem[5924] ;
wire \u_lsu.pmem[5925] ;
wire \u_lsu.pmem[5926] ;
wire \u_lsu.pmem[5927] ;
wire \u_lsu.pmem[5928] ;
wire \u_lsu.pmem[5929] ;
wire \u_lsu.pmem[5930] ;
wire \u_lsu.pmem[5931] ;
wire \u_lsu.pmem[5932] ;
wire \u_lsu.pmem[5933] ;
wire \u_lsu.pmem[5934] ;
wire \u_lsu.pmem[5935] ;
wire \u_lsu.pmem[5936] ;
wire \u_lsu.pmem[5937] ;
wire \u_lsu.pmem[5938] ;
wire \u_lsu.pmem[5939] ;
wire \u_lsu.pmem[5940] ;
wire \u_lsu.pmem[5941] ;
wire \u_lsu.pmem[5942] ;
wire \u_lsu.pmem[5943] ;
wire \u_lsu.pmem[5944] ;
wire \u_lsu.pmem[5945] ;
wire \u_lsu.pmem[5946] ;
wire \u_lsu.pmem[5947] ;
wire \u_lsu.pmem[5948] ;
wire \u_lsu.pmem[5949] ;
wire \u_lsu.pmem[5950] ;
wire \u_lsu.pmem[5951] ;
wire \u_lsu.pmem[5952] ;
wire \u_lsu.pmem[5953] ;
wire \u_lsu.pmem[5954] ;
wire \u_lsu.pmem[5955] ;
wire \u_lsu.pmem[5956] ;
wire \u_lsu.pmem[5957] ;
wire \u_lsu.pmem[5958] ;
wire \u_lsu.pmem[5959] ;
wire \u_lsu.pmem[5960] ;
wire \u_lsu.pmem[5961] ;
wire \u_lsu.pmem[5962] ;
wire \u_lsu.pmem[5963] ;
wire \u_lsu.pmem[5964] ;
wire \u_lsu.pmem[5965] ;
wire \u_lsu.pmem[5966] ;
wire \u_lsu.pmem[5967] ;
wire \u_lsu.pmem[5968] ;
wire \u_lsu.pmem[5969] ;
wire \u_lsu.pmem[5970] ;
wire \u_lsu.pmem[5971] ;
wire \u_lsu.pmem[5972] ;
wire \u_lsu.pmem[5973] ;
wire \u_lsu.pmem[5974] ;
wire \u_lsu.pmem[5975] ;
wire \u_lsu.pmem[5976] ;
wire \u_lsu.pmem[5977] ;
wire \u_lsu.pmem[5978] ;
wire \u_lsu.pmem[5979] ;
wire \u_lsu.pmem[5980] ;
wire \u_lsu.pmem[5981] ;
wire \u_lsu.pmem[5982] ;
wire \u_lsu.pmem[5983] ;
wire \u_lsu.pmem[5984] ;
wire \u_lsu.pmem[5985] ;
wire \u_lsu.pmem[5986] ;
wire \u_lsu.pmem[5987] ;
wire \u_lsu.pmem[5988] ;
wire \u_lsu.pmem[5989] ;
wire \u_lsu.pmem[5990] ;
wire \u_lsu.pmem[5991] ;
wire \u_lsu.pmem[5992] ;
wire \u_lsu.pmem[5993] ;
wire \u_lsu.pmem[5994] ;
wire \u_lsu.pmem[5995] ;
wire \u_lsu.pmem[5996] ;
wire \u_lsu.pmem[5997] ;
wire \u_lsu.pmem[5998] ;
wire \u_lsu.pmem[5999] ;
wire \u_lsu.pmem[6000] ;
wire \u_lsu.pmem[6001] ;
wire \u_lsu.pmem[6002] ;
wire \u_lsu.pmem[6003] ;
wire \u_lsu.pmem[6004] ;
wire \u_lsu.pmem[6005] ;
wire \u_lsu.pmem[6006] ;
wire \u_lsu.pmem[6007] ;
wire \u_lsu.pmem[6008] ;
wire \u_lsu.pmem[6009] ;
wire \u_lsu.pmem[6010] ;
wire \u_lsu.pmem[6011] ;
wire \u_lsu.pmem[6012] ;
wire \u_lsu.pmem[6013] ;
wire \u_lsu.pmem[6014] ;
wire \u_lsu.pmem[6015] ;
wire \u_lsu.pmem[6016] ;
wire \u_lsu.pmem[6017] ;
wire \u_lsu.pmem[6018] ;
wire \u_lsu.pmem[6019] ;
wire \u_lsu.pmem[6020] ;
wire \u_lsu.pmem[6021] ;
wire \u_lsu.pmem[6022] ;
wire \u_lsu.pmem[6023] ;
wire \u_lsu.pmem[6024] ;
wire \u_lsu.pmem[6025] ;
wire \u_lsu.pmem[6026] ;
wire \u_lsu.pmem[6027] ;
wire \u_lsu.pmem[6028] ;
wire \u_lsu.pmem[6029] ;
wire \u_lsu.pmem[6030] ;
wire \u_lsu.pmem[6031] ;
wire \u_lsu.pmem[6032] ;
wire \u_lsu.pmem[6033] ;
wire \u_lsu.pmem[6034] ;
wire \u_lsu.pmem[6035] ;
wire \u_lsu.pmem[6036] ;
wire \u_lsu.pmem[6037] ;
wire \u_lsu.pmem[6038] ;
wire \u_lsu.pmem[6039] ;
wire \u_lsu.pmem[6040] ;
wire \u_lsu.pmem[6041] ;
wire \u_lsu.pmem[6042] ;
wire \u_lsu.pmem[6043] ;
wire \u_lsu.pmem[6044] ;
wire \u_lsu.pmem[6045] ;
wire \u_lsu.pmem[6046] ;
wire \u_lsu.pmem[6047] ;
wire \u_lsu.pmem[6048] ;
wire \u_lsu.pmem[6049] ;
wire \u_lsu.pmem[6050] ;
wire \u_lsu.pmem[6051] ;
wire \u_lsu.pmem[6052] ;
wire \u_lsu.pmem[6053] ;
wire \u_lsu.pmem[6054] ;
wire \u_lsu.pmem[6055] ;
wire \u_lsu.pmem[6056] ;
wire \u_lsu.pmem[6057] ;
wire \u_lsu.pmem[6058] ;
wire \u_lsu.pmem[6059] ;
wire \u_lsu.pmem[6060] ;
wire \u_lsu.pmem[6061] ;
wire \u_lsu.pmem[6062] ;
wire \u_lsu.pmem[6063] ;
wire \u_lsu.pmem[6064] ;
wire \u_lsu.pmem[6065] ;
wire \u_lsu.pmem[6066] ;
wire \u_lsu.pmem[6067] ;
wire \u_lsu.pmem[6068] ;
wire \u_lsu.pmem[6069] ;
wire \u_lsu.pmem[6070] ;
wire \u_lsu.pmem[6071] ;
wire \u_lsu.pmem[6072] ;
wire \u_lsu.pmem[6073] ;
wire \u_lsu.pmem[6074] ;
wire \u_lsu.pmem[6075] ;
wire \u_lsu.pmem[6076] ;
wire \u_lsu.pmem[6077] ;
wire \u_lsu.pmem[6078] ;
wire \u_lsu.pmem[6079] ;
wire \u_lsu.pmem[6080] ;
wire \u_lsu.pmem[6081] ;
wire \u_lsu.pmem[6082] ;
wire \u_lsu.pmem[6083] ;
wire \u_lsu.pmem[6084] ;
wire \u_lsu.pmem[6085] ;
wire \u_lsu.pmem[6086] ;
wire \u_lsu.pmem[6087] ;
wire \u_lsu.pmem[6088] ;
wire \u_lsu.pmem[6089] ;
wire \u_lsu.pmem[6090] ;
wire \u_lsu.pmem[6091] ;
wire \u_lsu.pmem[6092] ;
wire \u_lsu.pmem[6093] ;
wire \u_lsu.pmem[6094] ;
wire \u_lsu.pmem[6095] ;
wire \u_lsu.pmem[6096] ;
wire \u_lsu.pmem[6097] ;
wire \u_lsu.pmem[6098] ;
wire \u_lsu.pmem[6099] ;
wire \u_lsu.pmem[6100] ;
wire \u_lsu.pmem[6101] ;
wire \u_lsu.pmem[6102] ;
wire \u_lsu.pmem[6103] ;
wire \u_lsu.pmem[6104] ;
wire \u_lsu.pmem[6105] ;
wire \u_lsu.pmem[6106] ;
wire \u_lsu.pmem[6107] ;
wire \u_lsu.pmem[6108] ;
wire \u_lsu.pmem[6109] ;
wire \u_lsu.pmem[6110] ;
wire \u_lsu.pmem[6111] ;
wire \u_lsu.pmem[6112] ;
wire \u_lsu.pmem[6113] ;
wire \u_lsu.pmem[6114] ;
wire \u_lsu.pmem[6115] ;
wire \u_lsu.pmem[6116] ;
wire \u_lsu.pmem[6117] ;
wire \u_lsu.pmem[6118] ;
wire \u_lsu.pmem[6119] ;
wire \u_lsu.pmem[6120] ;
wire \u_lsu.pmem[6121] ;
wire \u_lsu.pmem[6122] ;
wire \u_lsu.pmem[6123] ;
wire \u_lsu.pmem[6124] ;
wire \u_lsu.pmem[6125] ;
wire \u_lsu.pmem[6126] ;
wire \u_lsu.pmem[6127] ;
wire \u_lsu.pmem[6128] ;
wire \u_lsu.pmem[6129] ;
wire \u_lsu.pmem[6130] ;
wire \u_lsu.pmem[6131] ;
wire \u_lsu.pmem[6132] ;
wire \u_lsu.pmem[6133] ;
wire \u_lsu.pmem[6134] ;
wire \u_lsu.pmem[6135] ;
wire \u_lsu.pmem[6136] ;
wire \u_lsu.pmem[6137] ;
wire \u_lsu.pmem[6138] ;
wire \u_lsu.pmem[6139] ;
wire \u_lsu.pmem[6140] ;
wire \u_lsu.pmem[6141] ;
wire \u_lsu.pmem[6142] ;
wire \u_lsu.pmem[6143] ;
wire \u_lsu.pmem[6144] ;
wire \u_lsu.pmem[6145] ;
wire \u_lsu.pmem[6146] ;
wire \u_lsu.pmem[6147] ;
wire \u_lsu.pmem[6148] ;
wire \u_lsu.pmem[6149] ;
wire \u_lsu.pmem[6150] ;
wire \u_lsu.pmem[6151] ;
wire \u_lsu.pmem[6152] ;
wire \u_lsu.pmem[6153] ;
wire \u_lsu.pmem[6154] ;
wire \u_lsu.pmem[6155] ;
wire \u_lsu.pmem[6156] ;
wire \u_lsu.pmem[6157] ;
wire \u_lsu.pmem[6158] ;
wire \u_lsu.pmem[6159] ;
wire \u_lsu.pmem[6160] ;
wire \u_lsu.pmem[6161] ;
wire \u_lsu.pmem[6162] ;
wire \u_lsu.pmem[6163] ;
wire \u_lsu.pmem[6164] ;
wire \u_lsu.pmem[6165] ;
wire \u_lsu.pmem[6166] ;
wire \u_lsu.pmem[6167] ;
wire \u_lsu.pmem[6168] ;
wire \u_lsu.pmem[6169] ;
wire \u_lsu.pmem[6170] ;
wire \u_lsu.pmem[6171] ;
wire \u_lsu.pmem[6172] ;
wire \u_lsu.pmem[6173] ;
wire \u_lsu.pmem[6174] ;
wire \u_lsu.pmem[6175] ;
wire \u_lsu.pmem[6176] ;
wire \u_lsu.pmem[6177] ;
wire \u_lsu.pmem[6178] ;
wire \u_lsu.pmem[6179] ;
wire \u_lsu.pmem[6180] ;
wire \u_lsu.pmem[6181] ;
wire \u_lsu.pmem[6182] ;
wire \u_lsu.pmem[6183] ;
wire \u_lsu.pmem[6184] ;
wire \u_lsu.pmem[6185] ;
wire \u_lsu.pmem[6186] ;
wire \u_lsu.pmem[6187] ;
wire \u_lsu.pmem[6188] ;
wire \u_lsu.pmem[6189] ;
wire \u_lsu.pmem[6190] ;
wire \u_lsu.pmem[6191] ;
wire \u_lsu.pmem[6192] ;
wire \u_lsu.pmem[6193] ;
wire \u_lsu.pmem[6194] ;
wire \u_lsu.pmem[6195] ;
wire \u_lsu.pmem[6196] ;
wire \u_lsu.pmem[6197] ;
wire \u_lsu.pmem[6198] ;
wire \u_lsu.pmem[6199] ;
wire \u_lsu.pmem[6200] ;
wire \u_lsu.pmem[6201] ;
wire \u_lsu.pmem[6202] ;
wire \u_lsu.pmem[6203] ;
wire \u_lsu.pmem[6204] ;
wire \u_lsu.pmem[6205] ;
wire \u_lsu.pmem[6206] ;
wire \u_lsu.pmem[6207] ;
wire \u_lsu.pmem[6208] ;
wire \u_lsu.pmem[6209] ;
wire \u_lsu.pmem[6210] ;
wire \u_lsu.pmem[6211] ;
wire \u_lsu.pmem[6212] ;
wire \u_lsu.pmem[6213] ;
wire \u_lsu.pmem[6214] ;
wire \u_lsu.pmem[6215] ;
wire \u_lsu.pmem[6216] ;
wire \u_lsu.pmem[6217] ;
wire \u_lsu.pmem[6218] ;
wire \u_lsu.pmem[6219] ;
wire \u_lsu.pmem[6220] ;
wire \u_lsu.pmem[6221] ;
wire \u_lsu.pmem[6222] ;
wire \u_lsu.pmem[6223] ;
wire \u_lsu.pmem[6224] ;
wire \u_lsu.pmem[6225] ;
wire \u_lsu.pmem[6226] ;
wire \u_lsu.pmem[6227] ;
wire \u_lsu.pmem[6228] ;
wire \u_lsu.pmem[6229] ;
wire \u_lsu.pmem[6230] ;
wire \u_lsu.pmem[6231] ;
wire \u_lsu.pmem[6232] ;
wire \u_lsu.pmem[6233] ;
wire \u_lsu.pmem[6234] ;
wire \u_lsu.pmem[6235] ;
wire \u_lsu.pmem[6236] ;
wire \u_lsu.pmem[6237] ;
wire \u_lsu.pmem[6238] ;
wire \u_lsu.pmem[6239] ;
wire \u_lsu.pmem[6240] ;
wire \u_lsu.pmem[6241] ;
wire \u_lsu.pmem[6242] ;
wire \u_lsu.pmem[6243] ;
wire \u_lsu.pmem[6244] ;
wire \u_lsu.pmem[6245] ;
wire \u_lsu.pmem[6246] ;
wire \u_lsu.pmem[6247] ;
wire \u_lsu.pmem[6248] ;
wire \u_lsu.pmem[6249] ;
wire \u_lsu.pmem[6250] ;
wire \u_lsu.pmem[6251] ;
wire \u_lsu.pmem[6252] ;
wire \u_lsu.pmem[6253] ;
wire \u_lsu.pmem[6254] ;
wire \u_lsu.pmem[6255] ;
wire \u_lsu.pmem[6256] ;
wire \u_lsu.pmem[6257] ;
wire \u_lsu.pmem[6258] ;
wire \u_lsu.pmem[6259] ;
wire \u_lsu.pmem[6260] ;
wire \u_lsu.pmem[6261] ;
wire \u_lsu.pmem[6262] ;
wire \u_lsu.pmem[6263] ;
wire \u_lsu.pmem[6264] ;
wire \u_lsu.pmem[6265] ;
wire \u_lsu.pmem[6266] ;
wire \u_lsu.pmem[6267] ;
wire \u_lsu.pmem[6268] ;
wire \u_lsu.pmem[6269] ;
wire \u_lsu.pmem[6270] ;
wire \u_lsu.pmem[6271] ;
wire \u_lsu.pmem[6272] ;
wire \u_lsu.pmem[6273] ;
wire \u_lsu.pmem[6274] ;
wire \u_lsu.pmem[6275] ;
wire \u_lsu.pmem[6276] ;
wire \u_lsu.pmem[6277] ;
wire \u_lsu.pmem[6278] ;
wire \u_lsu.pmem[6279] ;
wire \u_lsu.pmem[6280] ;
wire \u_lsu.pmem[6281] ;
wire \u_lsu.pmem[6282] ;
wire \u_lsu.pmem[6283] ;
wire \u_lsu.pmem[6284] ;
wire \u_lsu.pmem[6285] ;
wire \u_lsu.pmem[6286] ;
wire \u_lsu.pmem[6287] ;
wire \u_lsu.pmem[6288] ;
wire \u_lsu.pmem[6289] ;
wire \u_lsu.pmem[6290] ;
wire \u_lsu.pmem[6291] ;
wire \u_lsu.pmem[6292] ;
wire \u_lsu.pmem[6293] ;
wire \u_lsu.pmem[6294] ;
wire \u_lsu.pmem[6295] ;
wire \u_lsu.pmem[6296] ;
wire \u_lsu.pmem[6297] ;
wire \u_lsu.pmem[6298] ;
wire \u_lsu.pmem[6299] ;
wire \u_lsu.pmem[6300] ;
wire \u_lsu.pmem[6301] ;
wire \u_lsu.pmem[6302] ;
wire \u_lsu.pmem[6303] ;
wire \u_lsu.pmem[6304] ;
wire \u_lsu.pmem[6305] ;
wire \u_lsu.pmem[6306] ;
wire \u_lsu.pmem[6307] ;
wire \u_lsu.pmem[6308] ;
wire \u_lsu.pmem[6309] ;
wire \u_lsu.pmem[6310] ;
wire \u_lsu.pmem[6311] ;
wire \u_lsu.pmem[6312] ;
wire \u_lsu.pmem[6313] ;
wire \u_lsu.pmem[6314] ;
wire \u_lsu.pmem[6315] ;
wire \u_lsu.pmem[6316] ;
wire \u_lsu.pmem[6317] ;
wire \u_lsu.pmem[6318] ;
wire \u_lsu.pmem[6319] ;
wire \u_lsu.pmem[6320] ;
wire \u_lsu.pmem[6321] ;
wire \u_lsu.pmem[6322] ;
wire \u_lsu.pmem[6323] ;
wire \u_lsu.pmem[6324] ;
wire \u_lsu.pmem[6325] ;
wire \u_lsu.pmem[6326] ;
wire \u_lsu.pmem[6327] ;
wire \u_lsu.pmem[6328] ;
wire \u_lsu.pmem[6329] ;
wire \u_lsu.pmem[6330] ;
wire \u_lsu.pmem[6331] ;
wire \u_lsu.pmem[6332] ;
wire \u_lsu.pmem[6333] ;
wire \u_lsu.pmem[6334] ;
wire \u_lsu.pmem[6335] ;
wire \u_lsu.pmem[6336] ;
wire \u_lsu.pmem[6337] ;
wire \u_lsu.pmem[6338] ;
wire \u_lsu.pmem[6339] ;
wire \u_lsu.pmem[6340] ;
wire \u_lsu.pmem[6341] ;
wire \u_lsu.pmem[6342] ;
wire \u_lsu.pmem[6343] ;
wire \u_lsu.pmem[6344] ;
wire \u_lsu.pmem[6345] ;
wire \u_lsu.pmem[6346] ;
wire \u_lsu.pmem[6347] ;
wire \u_lsu.pmem[6348] ;
wire \u_lsu.pmem[6349] ;
wire \u_lsu.pmem[6350] ;
wire \u_lsu.pmem[6351] ;
wire \u_lsu.pmem[6352] ;
wire \u_lsu.pmem[6353] ;
wire \u_lsu.pmem[6354] ;
wire \u_lsu.pmem[6355] ;
wire \u_lsu.pmem[6356] ;
wire \u_lsu.pmem[6357] ;
wire \u_lsu.pmem[6358] ;
wire \u_lsu.pmem[6359] ;
wire \u_lsu.pmem[6360] ;
wire \u_lsu.pmem[6361] ;
wire \u_lsu.pmem[6362] ;
wire \u_lsu.pmem[6363] ;
wire \u_lsu.pmem[6364] ;
wire \u_lsu.pmem[6365] ;
wire \u_lsu.pmem[6366] ;
wire \u_lsu.pmem[6367] ;
wire \u_lsu.pmem[6368] ;
wire \u_lsu.pmem[6369] ;
wire \u_lsu.pmem[6370] ;
wire \u_lsu.pmem[6371] ;
wire \u_lsu.pmem[6372] ;
wire \u_lsu.pmem[6373] ;
wire \u_lsu.pmem[6374] ;
wire \u_lsu.pmem[6375] ;
wire \u_lsu.pmem[6376] ;
wire \u_lsu.pmem[6377] ;
wire \u_lsu.pmem[6378] ;
wire \u_lsu.pmem[6379] ;
wire \u_lsu.pmem[6380] ;
wire \u_lsu.pmem[6381] ;
wire \u_lsu.pmem[6382] ;
wire \u_lsu.pmem[6383] ;
wire \u_lsu.pmem[6384] ;
wire \u_lsu.pmem[6385] ;
wire \u_lsu.pmem[6386] ;
wire \u_lsu.pmem[6387] ;
wire \u_lsu.pmem[6388] ;
wire \u_lsu.pmem[6389] ;
wire \u_lsu.pmem[6390] ;
wire \u_lsu.pmem[6391] ;
wire \u_lsu.pmem[6392] ;
wire \u_lsu.pmem[6393] ;
wire \u_lsu.pmem[6394] ;
wire \u_lsu.pmem[6395] ;
wire \u_lsu.pmem[6396] ;
wire \u_lsu.pmem[6397] ;
wire \u_lsu.pmem[6398] ;
wire \u_lsu.pmem[6399] ;
wire \u_lsu.pmem[6400] ;
wire \u_lsu.pmem[6401] ;
wire \u_lsu.pmem[6402] ;
wire \u_lsu.pmem[6403] ;
wire \u_lsu.pmem[6404] ;
wire \u_lsu.pmem[6405] ;
wire \u_lsu.pmem[6406] ;
wire \u_lsu.pmem[6407] ;
wire \u_lsu.pmem[6408] ;
wire \u_lsu.pmem[6409] ;
wire \u_lsu.pmem[6410] ;
wire \u_lsu.pmem[6411] ;
wire \u_lsu.pmem[6412] ;
wire \u_lsu.pmem[6413] ;
wire \u_lsu.pmem[6414] ;
wire \u_lsu.pmem[6415] ;
wire \u_lsu.pmem[6416] ;
wire \u_lsu.pmem[6417] ;
wire \u_lsu.pmem[6418] ;
wire \u_lsu.pmem[6419] ;
wire \u_lsu.pmem[6420] ;
wire \u_lsu.pmem[6421] ;
wire \u_lsu.pmem[6422] ;
wire \u_lsu.pmem[6423] ;
wire \u_lsu.pmem[6424] ;
wire \u_lsu.pmem[6425] ;
wire \u_lsu.pmem[6426] ;
wire \u_lsu.pmem[6427] ;
wire \u_lsu.pmem[6428] ;
wire \u_lsu.pmem[6429] ;
wire \u_lsu.pmem[6430] ;
wire \u_lsu.pmem[6431] ;
wire \u_lsu.pmem[6432] ;
wire \u_lsu.pmem[6433] ;
wire \u_lsu.pmem[6434] ;
wire \u_lsu.pmem[6435] ;
wire \u_lsu.pmem[6436] ;
wire \u_lsu.pmem[6437] ;
wire \u_lsu.pmem[6438] ;
wire \u_lsu.pmem[6439] ;
wire \u_lsu.pmem[6440] ;
wire \u_lsu.pmem[6441] ;
wire \u_lsu.pmem[6442] ;
wire \u_lsu.pmem[6443] ;
wire \u_lsu.pmem[6444] ;
wire \u_lsu.pmem[6445] ;
wire \u_lsu.pmem[6446] ;
wire \u_lsu.pmem[6447] ;
wire \u_lsu.pmem[6448] ;
wire \u_lsu.pmem[6449] ;
wire \u_lsu.pmem[6450] ;
wire \u_lsu.pmem[6451] ;
wire \u_lsu.pmem[6452] ;
wire \u_lsu.pmem[6453] ;
wire \u_lsu.pmem[6454] ;
wire \u_lsu.pmem[6455] ;
wire \u_lsu.pmem[6456] ;
wire \u_lsu.pmem[6457] ;
wire \u_lsu.pmem[6458] ;
wire \u_lsu.pmem[6459] ;
wire \u_lsu.pmem[6460] ;
wire \u_lsu.pmem[6461] ;
wire \u_lsu.pmem[6462] ;
wire \u_lsu.pmem[6463] ;
wire \u_lsu.pmem[6464] ;
wire \u_lsu.pmem[6465] ;
wire \u_lsu.pmem[6466] ;
wire \u_lsu.pmem[6467] ;
wire \u_lsu.pmem[6468] ;
wire \u_lsu.pmem[6469] ;
wire \u_lsu.pmem[6470] ;
wire \u_lsu.pmem[6471] ;
wire \u_lsu.pmem[6472] ;
wire \u_lsu.pmem[6473] ;
wire \u_lsu.pmem[6474] ;
wire \u_lsu.pmem[6475] ;
wire \u_lsu.pmem[6476] ;
wire \u_lsu.pmem[6477] ;
wire \u_lsu.pmem[6478] ;
wire \u_lsu.pmem[6479] ;
wire \u_lsu.pmem[6480] ;
wire \u_lsu.pmem[6481] ;
wire \u_lsu.pmem[6482] ;
wire \u_lsu.pmem[6483] ;
wire \u_lsu.pmem[6484] ;
wire \u_lsu.pmem[6485] ;
wire \u_lsu.pmem[6486] ;
wire \u_lsu.pmem[6487] ;
wire \u_lsu.pmem[6488] ;
wire \u_lsu.pmem[6489] ;
wire \u_lsu.pmem[6490] ;
wire \u_lsu.pmem[6491] ;
wire \u_lsu.pmem[6492] ;
wire \u_lsu.pmem[6493] ;
wire \u_lsu.pmem[6494] ;
wire \u_lsu.pmem[6495] ;
wire \u_lsu.pmem[6496] ;
wire \u_lsu.pmem[6497] ;
wire \u_lsu.pmem[6498] ;
wire \u_lsu.pmem[6499] ;
wire \u_lsu.pmem[6500] ;
wire \u_lsu.pmem[6501] ;
wire \u_lsu.pmem[6502] ;
wire \u_lsu.pmem[6503] ;
wire \u_lsu.pmem[6504] ;
wire \u_lsu.pmem[6505] ;
wire \u_lsu.pmem[6506] ;
wire \u_lsu.pmem[6507] ;
wire \u_lsu.pmem[6508] ;
wire \u_lsu.pmem[6509] ;
wire \u_lsu.pmem[6510] ;
wire \u_lsu.pmem[6511] ;
wire \u_lsu.pmem[6512] ;
wire \u_lsu.pmem[6513] ;
wire \u_lsu.pmem[6514] ;
wire \u_lsu.pmem[6515] ;
wire \u_lsu.pmem[6516] ;
wire \u_lsu.pmem[6517] ;
wire \u_lsu.pmem[6518] ;
wire \u_lsu.pmem[6519] ;
wire \u_lsu.pmem[6520] ;
wire \u_lsu.pmem[6521] ;
wire \u_lsu.pmem[6522] ;
wire \u_lsu.pmem[6523] ;
wire \u_lsu.pmem[6524] ;
wire \u_lsu.pmem[6525] ;
wire \u_lsu.pmem[6526] ;
wire \u_lsu.pmem[6527] ;
wire \u_lsu.pmem[6528] ;
wire \u_lsu.pmem[6529] ;
wire \u_lsu.pmem[6530] ;
wire \u_lsu.pmem[6531] ;
wire \u_lsu.pmem[6532] ;
wire \u_lsu.pmem[6533] ;
wire \u_lsu.pmem[6534] ;
wire \u_lsu.pmem[6535] ;
wire \u_lsu.pmem[6536] ;
wire \u_lsu.pmem[6537] ;
wire \u_lsu.pmem[6538] ;
wire \u_lsu.pmem[6539] ;
wire \u_lsu.pmem[6540] ;
wire \u_lsu.pmem[6541] ;
wire \u_lsu.pmem[6542] ;
wire \u_lsu.pmem[6543] ;
wire \u_lsu.pmem[6544] ;
wire \u_lsu.pmem[6545] ;
wire \u_lsu.pmem[6546] ;
wire \u_lsu.pmem[6547] ;
wire \u_lsu.pmem[6548] ;
wire \u_lsu.pmem[6549] ;
wire \u_lsu.pmem[6550] ;
wire \u_lsu.pmem[6551] ;
wire \u_lsu.pmem[6552] ;
wire \u_lsu.pmem[6553] ;
wire \u_lsu.pmem[6554] ;
wire \u_lsu.pmem[6555] ;
wire \u_lsu.pmem[6556] ;
wire \u_lsu.pmem[6557] ;
wire \u_lsu.pmem[6558] ;
wire \u_lsu.pmem[6559] ;
wire \u_lsu.pmem[6560] ;
wire \u_lsu.pmem[6561] ;
wire \u_lsu.pmem[6562] ;
wire \u_lsu.pmem[6563] ;
wire \u_lsu.pmem[6564] ;
wire \u_lsu.pmem[6565] ;
wire \u_lsu.pmem[6566] ;
wire \u_lsu.pmem[6567] ;
wire \u_lsu.pmem[6568] ;
wire \u_lsu.pmem[6569] ;
wire \u_lsu.pmem[6570] ;
wire \u_lsu.pmem[6571] ;
wire \u_lsu.pmem[6572] ;
wire \u_lsu.pmem[6573] ;
wire \u_lsu.pmem[6574] ;
wire \u_lsu.pmem[6575] ;
wire \u_lsu.pmem[6576] ;
wire \u_lsu.pmem[6577] ;
wire \u_lsu.pmem[6578] ;
wire \u_lsu.pmem[6579] ;
wire \u_lsu.pmem[6580] ;
wire \u_lsu.pmem[6581] ;
wire \u_lsu.pmem[6582] ;
wire \u_lsu.pmem[6583] ;
wire \u_lsu.pmem[6584] ;
wire \u_lsu.pmem[6585] ;
wire \u_lsu.pmem[6586] ;
wire \u_lsu.pmem[6587] ;
wire \u_lsu.pmem[6588] ;
wire \u_lsu.pmem[6589] ;
wire \u_lsu.pmem[6590] ;
wire \u_lsu.pmem[6591] ;
wire \u_lsu.pmem[6592] ;
wire \u_lsu.pmem[6593] ;
wire \u_lsu.pmem[6594] ;
wire \u_lsu.pmem[6595] ;
wire \u_lsu.pmem[6596] ;
wire \u_lsu.pmem[6597] ;
wire \u_lsu.pmem[6598] ;
wire \u_lsu.pmem[6599] ;
wire \u_lsu.pmem[6600] ;
wire \u_lsu.pmem[6601] ;
wire \u_lsu.pmem[6602] ;
wire \u_lsu.pmem[6603] ;
wire \u_lsu.pmem[6604] ;
wire \u_lsu.pmem[6605] ;
wire \u_lsu.pmem[6606] ;
wire \u_lsu.pmem[6607] ;
wire \u_lsu.pmem[6608] ;
wire \u_lsu.pmem[6609] ;
wire \u_lsu.pmem[6610] ;
wire \u_lsu.pmem[6611] ;
wire \u_lsu.pmem[6612] ;
wire \u_lsu.pmem[6613] ;
wire \u_lsu.pmem[6614] ;
wire \u_lsu.pmem[6615] ;
wire \u_lsu.pmem[6616] ;
wire \u_lsu.pmem[6617] ;
wire \u_lsu.pmem[6618] ;
wire \u_lsu.pmem[6619] ;
wire \u_lsu.pmem[6620] ;
wire \u_lsu.pmem[6621] ;
wire \u_lsu.pmem[6622] ;
wire \u_lsu.pmem[6623] ;
wire \u_lsu.pmem[6624] ;
wire \u_lsu.pmem[6625] ;
wire \u_lsu.pmem[6626] ;
wire \u_lsu.pmem[6627] ;
wire \u_lsu.pmem[6628] ;
wire \u_lsu.pmem[6629] ;
wire \u_lsu.pmem[6630] ;
wire \u_lsu.pmem[6631] ;
wire \u_lsu.pmem[6632] ;
wire \u_lsu.pmem[6633] ;
wire \u_lsu.pmem[6634] ;
wire \u_lsu.pmem[6635] ;
wire \u_lsu.pmem[6636] ;
wire \u_lsu.pmem[6637] ;
wire \u_lsu.pmem[6638] ;
wire \u_lsu.pmem[6639] ;
wire \u_lsu.pmem[6640] ;
wire \u_lsu.pmem[6641] ;
wire \u_lsu.pmem[6642] ;
wire \u_lsu.pmem[6643] ;
wire \u_lsu.pmem[6644] ;
wire \u_lsu.pmem[6645] ;
wire \u_lsu.pmem[6646] ;
wire \u_lsu.pmem[6647] ;
wire \u_lsu.pmem[6648] ;
wire \u_lsu.pmem[6649] ;
wire \u_lsu.pmem[6650] ;
wire \u_lsu.pmem[6651] ;
wire \u_lsu.pmem[6652] ;
wire \u_lsu.pmem[6653] ;
wire \u_lsu.pmem[6654] ;
wire \u_lsu.pmem[6655] ;
wire \u_lsu.pmem[6656] ;
wire \u_lsu.pmem[6657] ;
wire \u_lsu.pmem[6658] ;
wire \u_lsu.pmem[6659] ;
wire \u_lsu.pmem[6660] ;
wire \u_lsu.pmem[6661] ;
wire \u_lsu.pmem[6662] ;
wire \u_lsu.pmem[6663] ;
wire \u_lsu.pmem[6664] ;
wire \u_lsu.pmem[6665] ;
wire \u_lsu.pmem[6666] ;
wire \u_lsu.pmem[6667] ;
wire \u_lsu.pmem[6668] ;
wire \u_lsu.pmem[6669] ;
wire \u_lsu.pmem[6670] ;
wire \u_lsu.pmem[6671] ;
wire \u_lsu.pmem[6672] ;
wire \u_lsu.pmem[6673] ;
wire \u_lsu.pmem[6674] ;
wire \u_lsu.pmem[6675] ;
wire \u_lsu.pmem[6676] ;
wire \u_lsu.pmem[6677] ;
wire \u_lsu.pmem[6678] ;
wire \u_lsu.pmem[6679] ;
wire \u_lsu.pmem[6680] ;
wire \u_lsu.pmem[6681] ;
wire \u_lsu.pmem[6682] ;
wire \u_lsu.pmem[6683] ;
wire \u_lsu.pmem[6684] ;
wire \u_lsu.pmem[6685] ;
wire \u_lsu.pmem[6686] ;
wire \u_lsu.pmem[6687] ;
wire \u_lsu.pmem[6688] ;
wire \u_lsu.pmem[6689] ;
wire \u_lsu.pmem[6690] ;
wire \u_lsu.pmem[6691] ;
wire \u_lsu.pmem[6692] ;
wire \u_lsu.pmem[6693] ;
wire \u_lsu.pmem[6694] ;
wire \u_lsu.pmem[6695] ;
wire \u_lsu.pmem[6696] ;
wire \u_lsu.pmem[6697] ;
wire \u_lsu.pmem[6698] ;
wire \u_lsu.pmem[6699] ;
wire \u_lsu.pmem[6700] ;
wire \u_lsu.pmem[6701] ;
wire \u_lsu.pmem[6702] ;
wire \u_lsu.pmem[6703] ;
wire \u_lsu.pmem[6704] ;
wire \u_lsu.pmem[6705] ;
wire \u_lsu.pmem[6706] ;
wire \u_lsu.pmem[6707] ;
wire \u_lsu.pmem[6708] ;
wire \u_lsu.pmem[6709] ;
wire \u_lsu.pmem[6710] ;
wire \u_lsu.pmem[6711] ;
wire \u_lsu.pmem[6712] ;
wire \u_lsu.pmem[6713] ;
wire \u_lsu.pmem[6714] ;
wire \u_lsu.pmem[6715] ;
wire \u_lsu.pmem[6716] ;
wire \u_lsu.pmem[6717] ;
wire \u_lsu.pmem[6718] ;
wire \u_lsu.pmem[6719] ;
wire \u_lsu.pmem[6720] ;
wire \u_lsu.pmem[6721] ;
wire \u_lsu.pmem[6722] ;
wire \u_lsu.pmem[6723] ;
wire \u_lsu.pmem[6724] ;
wire \u_lsu.pmem[6725] ;
wire \u_lsu.pmem[6726] ;
wire \u_lsu.pmem[6727] ;
wire \u_lsu.pmem[6728] ;
wire \u_lsu.pmem[6729] ;
wire \u_lsu.pmem[6730] ;
wire \u_lsu.pmem[6731] ;
wire \u_lsu.pmem[6732] ;
wire \u_lsu.pmem[6733] ;
wire \u_lsu.pmem[6734] ;
wire \u_lsu.pmem[6735] ;
wire \u_lsu.pmem[6736] ;
wire \u_lsu.pmem[6737] ;
wire \u_lsu.pmem[6738] ;
wire \u_lsu.pmem[6739] ;
wire \u_lsu.pmem[6740] ;
wire \u_lsu.pmem[6741] ;
wire \u_lsu.pmem[6742] ;
wire \u_lsu.pmem[6743] ;
wire \u_lsu.pmem[6744] ;
wire \u_lsu.pmem[6745] ;
wire \u_lsu.pmem[6746] ;
wire \u_lsu.pmem[6747] ;
wire \u_lsu.pmem[6748] ;
wire \u_lsu.pmem[6749] ;
wire \u_lsu.pmem[6750] ;
wire \u_lsu.pmem[6751] ;
wire \u_lsu.pmem[6752] ;
wire \u_lsu.pmem[6753] ;
wire \u_lsu.pmem[6754] ;
wire \u_lsu.pmem[6755] ;
wire \u_lsu.pmem[6756] ;
wire \u_lsu.pmem[6757] ;
wire \u_lsu.pmem[6758] ;
wire \u_lsu.pmem[6759] ;
wire \u_lsu.pmem[6760] ;
wire \u_lsu.pmem[6761] ;
wire \u_lsu.pmem[6762] ;
wire \u_lsu.pmem[6763] ;
wire \u_lsu.pmem[6764] ;
wire \u_lsu.pmem[6765] ;
wire \u_lsu.pmem[6766] ;
wire \u_lsu.pmem[6767] ;
wire \u_lsu.pmem[6768] ;
wire \u_lsu.pmem[6769] ;
wire \u_lsu.pmem[6770] ;
wire \u_lsu.pmem[6771] ;
wire \u_lsu.pmem[6772] ;
wire \u_lsu.pmem[6773] ;
wire \u_lsu.pmem[6774] ;
wire \u_lsu.pmem[6775] ;
wire \u_lsu.pmem[6776] ;
wire \u_lsu.pmem[6777] ;
wire \u_lsu.pmem[6778] ;
wire \u_lsu.pmem[6779] ;
wire \u_lsu.pmem[6780] ;
wire \u_lsu.pmem[6781] ;
wire \u_lsu.pmem[6782] ;
wire \u_lsu.pmem[6783] ;
wire \u_lsu.pmem[6784] ;
wire \u_lsu.pmem[6785] ;
wire \u_lsu.pmem[6786] ;
wire \u_lsu.pmem[6787] ;
wire \u_lsu.pmem[6788] ;
wire \u_lsu.pmem[6789] ;
wire \u_lsu.pmem[6790] ;
wire \u_lsu.pmem[6791] ;
wire \u_lsu.pmem[6792] ;
wire \u_lsu.pmem[6793] ;
wire \u_lsu.pmem[6794] ;
wire \u_lsu.pmem[6795] ;
wire \u_lsu.pmem[6796] ;
wire \u_lsu.pmem[6797] ;
wire \u_lsu.pmem[6798] ;
wire \u_lsu.pmem[6799] ;
wire \u_lsu.pmem[6800] ;
wire \u_lsu.pmem[6801] ;
wire \u_lsu.pmem[6802] ;
wire \u_lsu.pmem[6803] ;
wire \u_lsu.pmem[6804] ;
wire \u_lsu.pmem[6805] ;
wire \u_lsu.pmem[6806] ;
wire \u_lsu.pmem[6807] ;
wire \u_lsu.pmem[6808] ;
wire \u_lsu.pmem[6809] ;
wire \u_lsu.pmem[6810] ;
wire \u_lsu.pmem[6811] ;
wire \u_lsu.pmem[6812] ;
wire \u_lsu.pmem[6813] ;
wire \u_lsu.pmem[6814] ;
wire \u_lsu.pmem[6815] ;
wire \u_lsu.pmem[6816] ;
wire \u_lsu.pmem[6817] ;
wire \u_lsu.pmem[6818] ;
wire \u_lsu.pmem[6819] ;
wire \u_lsu.pmem[6820] ;
wire \u_lsu.pmem[6821] ;
wire \u_lsu.pmem[6822] ;
wire \u_lsu.pmem[6823] ;
wire \u_lsu.pmem[6824] ;
wire \u_lsu.pmem[6825] ;
wire \u_lsu.pmem[6826] ;
wire \u_lsu.pmem[6827] ;
wire \u_lsu.pmem[6828] ;
wire \u_lsu.pmem[6829] ;
wire \u_lsu.pmem[6830] ;
wire \u_lsu.pmem[6831] ;
wire \u_lsu.pmem[6832] ;
wire \u_lsu.pmem[6833] ;
wire \u_lsu.pmem[6834] ;
wire \u_lsu.pmem[6835] ;
wire \u_lsu.pmem[6836] ;
wire \u_lsu.pmem[6837] ;
wire \u_lsu.pmem[6838] ;
wire \u_lsu.pmem[6839] ;
wire \u_lsu.pmem[6840] ;
wire \u_lsu.pmem[6841] ;
wire \u_lsu.pmem[6842] ;
wire \u_lsu.pmem[6843] ;
wire \u_lsu.pmem[6844] ;
wire \u_lsu.pmem[6845] ;
wire \u_lsu.pmem[6846] ;
wire \u_lsu.pmem[6847] ;
wire \u_lsu.pmem[6848] ;
wire \u_lsu.pmem[6849] ;
wire \u_lsu.pmem[6850] ;
wire \u_lsu.pmem[6851] ;
wire \u_lsu.pmem[6852] ;
wire \u_lsu.pmem[6853] ;
wire \u_lsu.pmem[6854] ;
wire \u_lsu.pmem[6855] ;
wire \u_lsu.pmem[6856] ;
wire \u_lsu.pmem[6857] ;
wire \u_lsu.pmem[6858] ;
wire \u_lsu.pmem[6859] ;
wire \u_lsu.pmem[6860] ;
wire \u_lsu.pmem[6861] ;
wire \u_lsu.pmem[6862] ;
wire \u_lsu.pmem[6863] ;
wire \u_lsu.pmem[6864] ;
wire \u_lsu.pmem[6865] ;
wire \u_lsu.pmem[6866] ;
wire \u_lsu.pmem[6867] ;
wire \u_lsu.pmem[6868] ;
wire \u_lsu.pmem[6869] ;
wire \u_lsu.pmem[6870] ;
wire \u_lsu.pmem[6871] ;
wire \u_lsu.pmem[6872] ;
wire \u_lsu.pmem[6873] ;
wire \u_lsu.pmem[6874] ;
wire \u_lsu.pmem[6875] ;
wire \u_lsu.pmem[6876] ;
wire \u_lsu.pmem[6877] ;
wire \u_lsu.pmem[6878] ;
wire \u_lsu.pmem[6879] ;
wire \u_lsu.pmem[6880] ;
wire \u_lsu.pmem[6881] ;
wire \u_lsu.pmem[6882] ;
wire \u_lsu.pmem[6883] ;
wire \u_lsu.pmem[6884] ;
wire \u_lsu.pmem[6885] ;
wire \u_lsu.pmem[6886] ;
wire \u_lsu.pmem[6887] ;
wire \u_lsu.pmem[6888] ;
wire \u_lsu.pmem[6889] ;
wire \u_lsu.pmem[6890] ;
wire \u_lsu.pmem[6891] ;
wire \u_lsu.pmem[6892] ;
wire \u_lsu.pmem[6893] ;
wire \u_lsu.pmem[6894] ;
wire \u_lsu.pmem[6895] ;
wire \u_lsu.pmem[6896] ;
wire \u_lsu.pmem[6897] ;
wire \u_lsu.pmem[6898] ;
wire \u_lsu.pmem[6899] ;
wire \u_lsu.pmem[6900] ;
wire \u_lsu.pmem[6901] ;
wire \u_lsu.pmem[6902] ;
wire \u_lsu.pmem[6903] ;
wire \u_lsu.pmem[6904] ;
wire \u_lsu.pmem[6905] ;
wire \u_lsu.pmem[6906] ;
wire \u_lsu.pmem[6907] ;
wire \u_lsu.pmem[6908] ;
wire \u_lsu.pmem[6909] ;
wire \u_lsu.pmem[6910] ;
wire \u_lsu.pmem[6911] ;
wire \u_lsu.pmem[6912] ;
wire \u_lsu.pmem[6913] ;
wire \u_lsu.pmem[6914] ;
wire \u_lsu.pmem[6915] ;
wire \u_lsu.pmem[6916] ;
wire \u_lsu.pmem[6917] ;
wire \u_lsu.pmem[6918] ;
wire \u_lsu.pmem[6919] ;
wire \u_lsu.pmem[6920] ;
wire \u_lsu.pmem[6921] ;
wire \u_lsu.pmem[6922] ;
wire \u_lsu.pmem[6923] ;
wire \u_lsu.pmem[6924] ;
wire \u_lsu.pmem[6925] ;
wire \u_lsu.pmem[6926] ;
wire \u_lsu.pmem[6927] ;
wire \u_lsu.pmem[6928] ;
wire \u_lsu.pmem[6929] ;
wire \u_lsu.pmem[6930] ;
wire \u_lsu.pmem[6931] ;
wire \u_lsu.pmem[6932] ;
wire \u_lsu.pmem[6933] ;
wire \u_lsu.pmem[6934] ;
wire \u_lsu.pmem[6935] ;
wire \u_lsu.pmem[6936] ;
wire \u_lsu.pmem[6937] ;
wire \u_lsu.pmem[6938] ;
wire \u_lsu.pmem[6939] ;
wire \u_lsu.pmem[6940] ;
wire \u_lsu.pmem[6941] ;
wire \u_lsu.pmem[6942] ;
wire \u_lsu.pmem[6943] ;
wire \u_lsu.pmem[6944] ;
wire \u_lsu.pmem[6945] ;
wire \u_lsu.pmem[6946] ;
wire \u_lsu.pmem[6947] ;
wire \u_lsu.pmem[6948] ;
wire \u_lsu.pmem[6949] ;
wire \u_lsu.pmem[6950] ;
wire \u_lsu.pmem[6951] ;
wire \u_lsu.pmem[6952] ;
wire \u_lsu.pmem[6953] ;
wire \u_lsu.pmem[6954] ;
wire \u_lsu.pmem[6955] ;
wire \u_lsu.pmem[6956] ;
wire \u_lsu.pmem[6957] ;
wire \u_lsu.pmem[6958] ;
wire \u_lsu.pmem[6959] ;
wire \u_lsu.pmem[6960] ;
wire \u_lsu.pmem[6961] ;
wire \u_lsu.pmem[6962] ;
wire \u_lsu.pmem[6963] ;
wire \u_lsu.pmem[6964] ;
wire \u_lsu.pmem[6965] ;
wire \u_lsu.pmem[6966] ;
wire \u_lsu.pmem[6967] ;
wire \u_lsu.pmem[6968] ;
wire \u_lsu.pmem[6969] ;
wire \u_lsu.pmem[6970] ;
wire \u_lsu.pmem[6971] ;
wire \u_lsu.pmem[6972] ;
wire \u_lsu.pmem[6973] ;
wire \u_lsu.pmem[6974] ;
wire \u_lsu.pmem[6975] ;
wire \u_lsu.pmem[6976] ;
wire \u_lsu.pmem[6977] ;
wire \u_lsu.pmem[6978] ;
wire \u_lsu.pmem[6979] ;
wire \u_lsu.pmem[6980] ;
wire \u_lsu.pmem[6981] ;
wire \u_lsu.pmem[6982] ;
wire \u_lsu.pmem[6983] ;
wire \u_lsu.pmem[6984] ;
wire \u_lsu.pmem[6985] ;
wire \u_lsu.pmem[6986] ;
wire \u_lsu.pmem[6987] ;
wire \u_lsu.pmem[6988] ;
wire \u_lsu.pmem[6989] ;
wire \u_lsu.pmem[6990] ;
wire \u_lsu.pmem[6991] ;
wire \u_lsu.pmem[6992] ;
wire \u_lsu.pmem[6993] ;
wire \u_lsu.pmem[6994] ;
wire \u_lsu.pmem[6995] ;
wire \u_lsu.pmem[6996] ;
wire \u_lsu.pmem[6997] ;
wire \u_lsu.pmem[6998] ;
wire \u_lsu.pmem[6999] ;
wire \u_lsu.pmem[7000] ;
wire \u_lsu.pmem[7001] ;
wire \u_lsu.pmem[7002] ;
wire \u_lsu.pmem[7003] ;
wire \u_lsu.pmem[7004] ;
wire \u_lsu.pmem[7005] ;
wire \u_lsu.pmem[7006] ;
wire \u_lsu.pmem[7007] ;
wire \u_lsu.pmem[7008] ;
wire \u_lsu.pmem[7009] ;
wire \u_lsu.pmem[7010] ;
wire \u_lsu.pmem[7011] ;
wire \u_lsu.pmem[7012] ;
wire \u_lsu.pmem[7013] ;
wire \u_lsu.pmem[7014] ;
wire \u_lsu.pmem[7015] ;
wire \u_lsu.pmem[7016] ;
wire \u_lsu.pmem[7017] ;
wire \u_lsu.pmem[7018] ;
wire \u_lsu.pmem[7019] ;
wire \u_lsu.pmem[7020] ;
wire \u_lsu.pmem[7021] ;
wire \u_lsu.pmem[7022] ;
wire \u_lsu.pmem[7023] ;
wire \u_lsu.pmem[7024] ;
wire \u_lsu.pmem[7025] ;
wire \u_lsu.pmem[7026] ;
wire \u_lsu.pmem[7027] ;
wire \u_lsu.pmem[7028] ;
wire \u_lsu.pmem[7029] ;
wire \u_lsu.pmem[7030] ;
wire \u_lsu.pmem[7031] ;
wire \u_lsu.pmem[7032] ;
wire \u_lsu.pmem[7033] ;
wire \u_lsu.pmem[7034] ;
wire \u_lsu.pmem[7035] ;
wire \u_lsu.pmem[7036] ;
wire \u_lsu.pmem[7037] ;
wire \u_lsu.pmem[7038] ;
wire \u_lsu.pmem[7039] ;
wire \u_lsu.pmem[7040] ;
wire \u_lsu.pmem[7041] ;
wire \u_lsu.pmem[7042] ;
wire \u_lsu.pmem[7043] ;
wire \u_lsu.pmem[7044] ;
wire \u_lsu.pmem[7045] ;
wire \u_lsu.pmem[7046] ;
wire \u_lsu.pmem[7047] ;
wire \u_lsu.pmem[7048] ;
wire \u_lsu.pmem[7049] ;
wire \u_lsu.pmem[7050] ;
wire \u_lsu.pmem[7051] ;
wire \u_lsu.pmem[7052] ;
wire \u_lsu.pmem[7053] ;
wire \u_lsu.pmem[7054] ;
wire \u_lsu.pmem[7055] ;
wire \u_lsu.pmem[7056] ;
wire \u_lsu.pmem[7057] ;
wire \u_lsu.pmem[7058] ;
wire \u_lsu.pmem[7059] ;
wire \u_lsu.pmem[7060] ;
wire \u_lsu.pmem[7061] ;
wire \u_lsu.pmem[7062] ;
wire \u_lsu.pmem[7063] ;
wire \u_lsu.pmem[7064] ;
wire \u_lsu.pmem[7065] ;
wire \u_lsu.pmem[7066] ;
wire \u_lsu.pmem[7067] ;
wire \u_lsu.pmem[7068] ;
wire \u_lsu.pmem[7069] ;
wire \u_lsu.pmem[7070] ;
wire \u_lsu.pmem[7071] ;
wire \u_lsu.pmem[7072] ;
wire \u_lsu.pmem[7073] ;
wire \u_lsu.pmem[7074] ;
wire \u_lsu.pmem[7075] ;
wire \u_lsu.pmem[7076] ;
wire \u_lsu.pmem[7077] ;
wire \u_lsu.pmem[7078] ;
wire \u_lsu.pmem[7079] ;
wire \u_lsu.pmem[7080] ;
wire \u_lsu.pmem[7081] ;
wire \u_lsu.pmem[7082] ;
wire \u_lsu.pmem[7083] ;
wire \u_lsu.pmem[7084] ;
wire \u_lsu.pmem[7085] ;
wire \u_lsu.pmem[7086] ;
wire \u_lsu.pmem[7087] ;
wire \u_lsu.pmem[7088] ;
wire \u_lsu.pmem[7089] ;
wire \u_lsu.pmem[7090] ;
wire \u_lsu.pmem[7091] ;
wire \u_lsu.pmem[7092] ;
wire \u_lsu.pmem[7093] ;
wire \u_lsu.pmem[7094] ;
wire \u_lsu.pmem[7095] ;
wire \u_lsu.pmem[7096] ;
wire \u_lsu.pmem[7097] ;
wire \u_lsu.pmem[7098] ;
wire \u_lsu.pmem[7099] ;
wire \u_lsu.pmem[7100] ;
wire \u_lsu.pmem[7101] ;
wire \u_lsu.pmem[7102] ;
wire \u_lsu.pmem[7103] ;
wire \u_lsu.pmem[7104] ;
wire \u_lsu.pmem[7105] ;
wire \u_lsu.pmem[7106] ;
wire \u_lsu.pmem[7107] ;
wire \u_lsu.pmem[7108] ;
wire \u_lsu.pmem[7109] ;
wire \u_lsu.pmem[7110] ;
wire \u_lsu.pmem[7111] ;
wire \u_lsu.pmem[7112] ;
wire \u_lsu.pmem[7113] ;
wire \u_lsu.pmem[7114] ;
wire \u_lsu.pmem[7115] ;
wire \u_lsu.pmem[7116] ;
wire \u_lsu.pmem[7117] ;
wire \u_lsu.pmem[7118] ;
wire \u_lsu.pmem[7119] ;
wire \u_lsu.pmem[7120] ;
wire \u_lsu.pmem[7121] ;
wire \u_lsu.pmem[7122] ;
wire \u_lsu.pmem[7123] ;
wire \u_lsu.pmem[7124] ;
wire \u_lsu.pmem[7125] ;
wire \u_lsu.pmem[7126] ;
wire \u_lsu.pmem[7127] ;
wire \u_lsu.pmem[7128] ;
wire \u_lsu.pmem[7129] ;
wire \u_lsu.pmem[7130] ;
wire \u_lsu.pmem[7131] ;
wire \u_lsu.pmem[7132] ;
wire \u_lsu.pmem[7133] ;
wire \u_lsu.pmem[7134] ;
wire \u_lsu.pmem[7135] ;
wire \u_lsu.pmem[7136] ;
wire \u_lsu.pmem[7137] ;
wire \u_lsu.pmem[7138] ;
wire \u_lsu.pmem[7139] ;
wire \u_lsu.pmem[7140] ;
wire \u_lsu.pmem[7141] ;
wire \u_lsu.pmem[7142] ;
wire \u_lsu.pmem[7143] ;
wire \u_lsu.pmem[7144] ;
wire \u_lsu.pmem[7145] ;
wire \u_lsu.pmem[7146] ;
wire \u_lsu.pmem[7147] ;
wire \u_lsu.pmem[7148] ;
wire \u_lsu.pmem[7149] ;
wire \u_lsu.pmem[7150] ;
wire \u_lsu.pmem[7151] ;
wire \u_lsu.pmem[7152] ;
wire \u_lsu.pmem[7153] ;
wire \u_lsu.pmem[7154] ;
wire \u_lsu.pmem[7155] ;
wire \u_lsu.pmem[7156] ;
wire \u_lsu.pmem[7157] ;
wire \u_lsu.pmem[7158] ;
wire \u_lsu.pmem[7159] ;
wire \u_lsu.pmem[7160] ;
wire \u_lsu.pmem[7161] ;
wire \u_lsu.pmem[7162] ;
wire \u_lsu.pmem[7163] ;
wire \u_lsu.pmem[7164] ;
wire \u_lsu.pmem[7165] ;
wire \u_lsu.pmem[7166] ;
wire \u_lsu.pmem[7167] ;
wire \u_lsu.pmem[7168] ;
wire \u_lsu.pmem[7169] ;
wire \u_lsu.pmem[7170] ;
wire \u_lsu.pmem[7171] ;
wire \u_lsu.pmem[7172] ;
wire \u_lsu.pmem[7173] ;
wire \u_lsu.pmem[7174] ;
wire \u_lsu.pmem[7175] ;
wire \u_lsu.pmem[7176] ;
wire \u_lsu.pmem[7177] ;
wire \u_lsu.pmem[7178] ;
wire \u_lsu.pmem[7179] ;
wire \u_lsu.pmem[7180] ;
wire \u_lsu.pmem[7181] ;
wire \u_lsu.pmem[7182] ;
wire \u_lsu.pmem[7183] ;
wire \u_lsu.pmem[7184] ;
wire \u_lsu.pmem[7185] ;
wire \u_lsu.pmem[7186] ;
wire \u_lsu.pmem[7187] ;
wire \u_lsu.pmem[7188] ;
wire \u_lsu.pmem[7189] ;
wire \u_lsu.pmem[7190] ;
wire \u_lsu.pmem[7191] ;
wire \u_lsu.pmem[7192] ;
wire \u_lsu.pmem[7193] ;
wire \u_lsu.pmem[7194] ;
wire \u_lsu.pmem[7195] ;
wire \u_lsu.pmem[7196] ;
wire \u_lsu.pmem[7197] ;
wire \u_lsu.pmem[7198] ;
wire \u_lsu.pmem[7199] ;
wire \u_lsu.pmem[7200] ;
wire \u_lsu.pmem[7201] ;
wire \u_lsu.pmem[7202] ;
wire \u_lsu.pmem[7203] ;
wire \u_lsu.pmem[7204] ;
wire \u_lsu.pmem[7205] ;
wire \u_lsu.pmem[7206] ;
wire \u_lsu.pmem[7207] ;
wire \u_lsu.pmem[7208] ;
wire \u_lsu.pmem[7209] ;
wire \u_lsu.pmem[7210] ;
wire \u_lsu.pmem[7211] ;
wire \u_lsu.pmem[7212] ;
wire \u_lsu.pmem[7213] ;
wire \u_lsu.pmem[7214] ;
wire \u_lsu.pmem[7215] ;
wire \u_lsu.pmem[7216] ;
wire \u_lsu.pmem[7217] ;
wire \u_lsu.pmem[7218] ;
wire \u_lsu.pmem[7219] ;
wire \u_lsu.pmem[7220] ;
wire \u_lsu.pmem[7221] ;
wire \u_lsu.pmem[7222] ;
wire \u_lsu.pmem[7223] ;
wire \u_lsu.pmem[7224] ;
wire \u_lsu.pmem[7225] ;
wire \u_lsu.pmem[7226] ;
wire \u_lsu.pmem[7227] ;
wire \u_lsu.pmem[7228] ;
wire \u_lsu.pmem[7229] ;
wire \u_lsu.pmem[7230] ;
wire \u_lsu.pmem[7231] ;
wire \u_lsu.pmem[7232] ;
wire \u_lsu.pmem[7233] ;
wire \u_lsu.pmem[7234] ;
wire \u_lsu.pmem[7235] ;
wire \u_lsu.pmem[7236] ;
wire \u_lsu.pmem[7237] ;
wire \u_lsu.pmem[7238] ;
wire \u_lsu.pmem[7239] ;
wire \u_lsu.pmem[7240] ;
wire \u_lsu.pmem[7241] ;
wire \u_lsu.pmem[7242] ;
wire \u_lsu.pmem[7243] ;
wire \u_lsu.pmem[7244] ;
wire \u_lsu.pmem[7245] ;
wire \u_lsu.pmem[7246] ;
wire \u_lsu.pmem[7247] ;
wire \u_lsu.pmem[7248] ;
wire \u_lsu.pmem[7249] ;
wire \u_lsu.pmem[7250] ;
wire \u_lsu.pmem[7251] ;
wire \u_lsu.pmem[7252] ;
wire \u_lsu.pmem[7253] ;
wire \u_lsu.pmem[7254] ;
wire \u_lsu.pmem[7255] ;
wire \u_lsu.pmem[7256] ;
wire \u_lsu.pmem[7257] ;
wire \u_lsu.pmem[7258] ;
wire \u_lsu.pmem[7259] ;
wire \u_lsu.pmem[7260] ;
wire \u_lsu.pmem[7261] ;
wire \u_lsu.pmem[7262] ;
wire \u_lsu.pmem[7263] ;
wire \u_lsu.pmem[7264] ;
wire \u_lsu.pmem[7265] ;
wire \u_lsu.pmem[7266] ;
wire \u_lsu.pmem[7267] ;
wire \u_lsu.pmem[7268] ;
wire \u_lsu.pmem[7269] ;
wire \u_lsu.pmem[7270] ;
wire \u_lsu.pmem[7271] ;
wire \u_lsu.pmem[7272] ;
wire \u_lsu.pmem[7273] ;
wire \u_lsu.pmem[7274] ;
wire \u_lsu.pmem[7275] ;
wire \u_lsu.pmem[7276] ;
wire \u_lsu.pmem[7277] ;
wire \u_lsu.pmem[7278] ;
wire \u_lsu.pmem[7279] ;
wire \u_lsu.pmem[7280] ;
wire \u_lsu.pmem[7281] ;
wire \u_lsu.pmem[7282] ;
wire \u_lsu.pmem[7283] ;
wire \u_lsu.pmem[7284] ;
wire \u_lsu.pmem[7285] ;
wire \u_lsu.pmem[7286] ;
wire \u_lsu.pmem[7287] ;
wire \u_lsu.pmem[7288] ;
wire \u_lsu.pmem[7289] ;
wire \u_lsu.pmem[7290] ;
wire \u_lsu.pmem[7291] ;
wire \u_lsu.pmem[7292] ;
wire \u_lsu.pmem[7293] ;
wire \u_lsu.pmem[7294] ;
wire \u_lsu.pmem[7295] ;
wire \u_lsu.pmem[7296] ;
wire \u_lsu.pmem[7297] ;
wire \u_lsu.pmem[7298] ;
wire \u_lsu.pmem[7299] ;
wire \u_lsu.pmem[7300] ;
wire \u_lsu.pmem[7301] ;
wire \u_lsu.pmem[7302] ;
wire \u_lsu.pmem[7303] ;
wire \u_lsu.pmem[7304] ;
wire \u_lsu.pmem[7305] ;
wire \u_lsu.pmem[7306] ;
wire \u_lsu.pmem[7307] ;
wire \u_lsu.pmem[7308] ;
wire \u_lsu.pmem[7309] ;
wire \u_lsu.pmem[7310] ;
wire \u_lsu.pmem[7311] ;
wire \u_lsu.pmem[7312] ;
wire \u_lsu.pmem[7313] ;
wire \u_lsu.pmem[7314] ;
wire \u_lsu.pmem[7315] ;
wire \u_lsu.pmem[7316] ;
wire \u_lsu.pmem[7317] ;
wire \u_lsu.pmem[7318] ;
wire \u_lsu.pmem[7319] ;
wire \u_lsu.pmem[7320] ;
wire \u_lsu.pmem[7321] ;
wire \u_lsu.pmem[7322] ;
wire \u_lsu.pmem[7323] ;
wire \u_lsu.pmem[7324] ;
wire \u_lsu.pmem[7325] ;
wire \u_lsu.pmem[7326] ;
wire \u_lsu.pmem[7327] ;
wire \u_lsu.pmem[7328] ;
wire \u_lsu.pmem[7329] ;
wire \u_lsu.pmem[7330] ;
wire \u_lsu.pmem[7331] ;
wire \u_lsu.pmem[7332] ;
wire \u_lsu.pmem[7333] ;
wire \u_lsu.pmem[7334] ;
wire \u_lsu.pmem[7335] ;
wire \u_lsu.pmem[7336] ;
wire \u_lsu.pmem[7337] ;
wire \u_lsu.pmem[7338] ;
wire \u_lsu.pmem[7339] ;
wire \u_lsu.pmem[7340] ;
wire \u_lsu.pmem[7341] ;
wire \u_lsu.pmem[7342] ;
wire \u_lsu.pmem[7343] ;
wire \u_lsu.pmem[7344] ;
wire \u_lsu.pmem[7345] ;
wire \u_lsu.pmem[7346] ;
wire \u_lsu.pmem[7347] ;
wire \u_lsu.pmem[7348] ;
wire \u_lsu.pmem[7349] ;
wire \u_lsu.pmem[7350] ;
wire \u_lsu.pmem[7351] ;
wire \u_lsu.pmem[7352] ;
wire \u_lsu.pmem[7353] ;
wire \u_lsu.pmem[7354] ;
wire \u_lsu.pmem[7355] ;
wire \u_lsu.pmem[7356] ;
wire \u_lsu.pmem[7357] ;
wire \u_lsu.pmem[7358] ;
wire \u_lsu.pmem[7359] ;
wire \u_lsu.pmem[7360] ;
wire \u_lsu.pmem[7361] ;
wire \u_lsu.pmem[7362] ;
wire \u_lsu.pmem[7363] ;
wire \u_lsu.pmem[7364] ;
wire \u_lsu.pmem[7365] ;
wire \u_lsu.pmem[7366] ;
wire \u_lsu.pmem[7367] ;
wire \u_lsu.pmem[7368] ;
wire \u_lsu.pmem[7369] ;
wire \u_lsu.pmem[7370] ;
wire \u_lsu.pmem[7371] ;
wire \u_lsu.pmem[7372] ;
wire \u_lsu.pmem[7373] ;
wire \u_lsu.pmem[7374] ;
wire \u_lsu.pmem[7375] ;
wire \u_lsu.pmem[7376] ;
wire \u_lsu.pmem[7377] ;
wire \u_lsu.pmem[7378] ;
wire \u_lsu.pmem[7379] ;
wire \u_lsu.pmem[7380] ;
wire \u_lsu.pmem[7381] ;
wire \u_lsu.pmem[7382] ;
wire \u_lsu.pmem[7383] ;
wire \u_lsu.pmem[7384] ;
wire \u_lsu.pmem[7385] ;
wire \u_lsu.pmem[7386] ;
wire \u_lsu.pmem[7387] ;
wire \u_lsu.pmem[7388] ;
wire \u_lsu.pmem[7389] ;
wire \u_lsu.pmem[7390] ;
wire \u_lsu.pmem[7391] ;
wire \u_lsu.pmem[7392] ;
wire \u_lsu.pmem[7393] ;
wire \u_lsu.pmem[7394] ;
wire \u_lsu.pmem[7395] ;
wire \u_lsu.pmem[7396] ;
wire \u_lsu.pmem[7397] ;
wire \u_lsu.pmem[7398] ;
wire \u_lsu.pmem[7399] ;
wire \u_lsu.pmem[7400] ;
wire \u_lsu.pmem[7401] ;
wire \u_lsu.pmem[7402] ;
wire \u_lsu.pmem[7403] ;
wire \u_lsu.pmem[7404] ;
wire \u_lsu.pmem[7405] ;
wire \u_lsu.pmem[7406] ;
wire \u_lsu.pmem[7407] ;
wire \u_lsu.pmem[7408] ;
wire \u_lsu.pmem[7409] ;
wire \u_lsu.pmem[7410] ;
wire \u_lsu.pmem[7411] ;
wire \u_lsu.pmem[7412] ;
wire \u_lsu.pmem[7413] ;
wire \u_lsu.pmem[7414] ;
wire \u_lsu.pmem[7415] ;
wire \u_lsu.pmem[7416] ;
wire \u_lsu.pmem[7417] ;
wire \u_lsu.pmem[7418] ;
wire \u_lsu.pmem[7419] ;
wire \u_lsu.pmem[7420] ;
wire \u_lsu.pmem[7421] ;
wire \u_lsu.pmem[7422] ;
wire \u_lsu.pmem[7423] ;
wire \u_lsu.pmem[7424] ;
wire \u_lsu.pmem[7425] ;
wire \u_lsu.pmem[7426] ;
wire \u_lsu.pmem[7427] ;
wire \u_lsu.pmem[7428] ;
wire \u_lsu.pmem[7429] ;
wire \u_lsu.pmem[7430] ;
wire \u_lsu.pmem[7431] ;
wire \u_lsu.pmem[7432] ;
wire \u_lsu.pmem[7433] ;
wire \u_lsu.pmem[7434] ;
wire \u_lsu.pmem[7435] ;
wire \u_lsu.pmem[7436] ;
wire \u_lsu.pmem[7437] ;
wire \u_lsu.pmem[7438] ;
wire \u_lsu.pmem[7439] ;
wire \u_lsu.pmem[7440] ;
wire \u_lsu.pmem[7441] ;
wire \u_lsu.pmem[7442] ;
wire \u_lsu.pmem[7443] ;
wire \u_lsu.pmem[7444] ;
wire \u_lsu.pmem[7445] ;
wire \u_lsu.pmem[7446] ;
wire \u_lsu.pmem[7447] ;
wire \u_lsu.pmem[7448] ;
wire \u_lsu.pmem[7449] ;
wire \u_lsu.pmem[7450] ;
wire \u_lsu.pmem[7451] ;
wire \u_lsu.pmem[7452] ;
wire \u_lsu.pmem[7453] ;
wire \u_lsu.pmem[7454] ;
wire \u_lsu.pmem[7455] ;
wire \u_lsu.pmem[7456] ;
wire \u_lsu.pmem[7457] ;
wire \u_lsu.pmem[7458] ;
wire \u_lsu.pmem[7459] ;
wire \u_lsu.pmem[7460] ;
wire \u_lsu.pmem[7461] ;
wire \u_lsu.pmem[7462] ;
wire \u_lsu.pmem[7463] ;
wire \u_lsu.pmem[7464] ;
wire \u_lsu.pmem[7465] ;
wire \u_lsu.pmem[7466] ;
wire \u_lsu.pmem[7467] ;
wire \u_lsu.pmem[7468] ;
wire \u_lsu.pmem[7469] ;
wire \u_lsu.pmem[7470] ;
wire \u_lsu.pmem[7471] ;
wire \u_lsu.pmem[7472] ;
wire \u_lsu.pmem[7473] ;
wire \u_lsu.pmem[7474] ;
wire \u_lsu.pmem[7475] ;
wire \u_lsu.pmem[7476] ;
wire \u_lsu.pmem[7477] ;
wire \u_lsu.pmem[7478] ;
wire \u_lsu.pmem[7479] ;
wire \u_lsu.pmem[7480] ;
wire \u_lsu.pmem[7481] ;
wire \u_lsu.pmem[7482] ;
wire \u_lsu.pmem[7483] ;
wire \u_lsu.pmem[7484] ;
wire \u_lsu.pmem[7485] ;
wire \u_lsu.pmem[7486] ;
wire \u_lsu.pmem[7487] ;
wire \u_lsu.pmem[7488] ;
wire \u_lsu.pmem[7489] ;
wire \u_lsu.pmem[7490] ;
wire \u_lsu.pmem[7491] ;
wire \u_lsu.pmem[7492] ;
wire \u_lsu.pmem[7493] ;
wire \u_lsu.pmem[7494] ;
wire \u_lsu.pmem[7495] ;
wire \u_lsu.pmem[7496] ;
wire \u_lsu.pmem[7497] ;
wire \u_lsu.pmem[7498] ;
wire \u_lsu.pmem[7499] ;
wire \u_lsu.pmem[7500] ;
wire \u_lsu.pmem[7501] ;
wire \u_lsu.pmem[7502] ;
wire \u_lsu.pmem[7503] ;
wire \u_lsu.pmem[7504] ;
wire \u_lsu.pmem[7505] ;
wire \u_lsu.pmem[7506] ;
wire \u_lsu.pmem[7507] ;
wire \u_lsu.pmem[7508] ;
wire \u_lsu.pmem[7509] ;
wire \u_lsu.pmem[7510] ;
wire \u_lsu.pmem[7511] ;
wire \u_lsu.pmem[7512] ;
wire \u_lsu.pmem[7513] ;
wire \u_lsu.pmem[7514] ;
wire \u_lsu.pmem[7515] ;
wire \u_lsu.pmem[7516] ;
wire \u_lsu.pmem[7517] ;
wire \u_lsu.pmem[7518] ;
wire \u_lsu.pmem[7519] ;
wire \u_lsu.pmem[7520] ;
wire \u_lsu.pmem[7521] ;
wire \u_lsu.pmem[7522] ;
wire \u_lsu.pmem[7523] ;
wire \u_lsu.pmem[7524] ;
wire \u_lsu.pmem[7525] ;
wire \u_lsu.pmem[7526] ;
wire \u_lsu.pmem[7527] ;
wire \u_lsu.pmem[7528] ;
wire \u_lsu.pmem[7529] ;
wire \u_lsu.pmem[7530] ;
wire \u_lsu.pmem[7531] ;
wire \u_lsu.pmem[7532] ;
wire \u_lsu.pmem[7533] ;
wire \u_lsu.pmem[7534] ;
wire \u_lsu.pmem[7535] ;
wire \u_lsu.pmem[7536] ;
wire \u_lsu.pmem[7537] ;
wire \u_lsu.pmem[7538] ;
wire \u_lsu.pmem[7539] ;
wire \u_lsu.pmem[7540] ;
wire \u_lsu.pmem[7541] ;
wire \u_lsu.pmem[7542] ;
wire \u_lsu.pmem[7543] ;
wire \u_lsu.pmem[7544] ;
wire \u_lsu.pmem[7545] ;
wire \u_lsu.pmem[7546] ;
wire \u_lsu.pmem[7547] ;
wire \u_lsu.pmem[7548] ;
wire \u_lsu.pmem[7549] ;
wire \u_lsu.pmem[7550] ;
wire \u_lsu.pmem[7551] ;
wire \u_lsu.pmem[7552] ;
wire \u_lsu.pmem[7553] ;
wire \u_lsu.pmem[7554] ;
wire \u_lsu.pmem[7555] ;
wire \u_lsu.pmem[7556] ;
wire \u_lsu.pmem[7557] ;
wire \u_lsu.pmem[7558] ;
wire \u_lsu.pmem[7559] ;
wire \u_lsu.pmem[7560] ;
wire \u_lsu.pmem[7561] ;
wire \u_lsu.pmem[7562] ;
wire \u_lsu.pmem[7563] ;
wire \u_lsu.pmem[7564] ;
wire \u_lsu.pmem[7565] ;
wire \u_lsu.pmem[7566] ;
wire \u_lsu.pmem[7567] ;
wire \u_lsu.pmem[7568] ;
wire \u_lsu.pmem[7569] ;
wire \u_lsu.pmem[7570] ;
wire \u_lsu.pmem[7571] ;
wire \u_lsu.pmem[7572] ;
wire \u_lsu.pmem[7573] ;
wire \u_lsu.pmem[7574] ;
wire \u_lsu.pmem[7575] ;
wire \u_lsu.pmem[7576] ;
wire \u_lsu.pmem[7577] ;
wire \u_lsu.pmem[7578] ;
wire \u_lsu.pmem[7579] ;
wire \u_lsu.pmem[7580] ;
wire \u_lsu.pmem[7581] ;
wire \u_lsu.pmem[7582] ;
wire \u_lsu.pmem[7583] ;
wire \u_lsu.pmem[7584] ;
wire \u_lsu.pmem[7585] ;
wire \u_lsu.pmem[7586] ;
wire \u_lsu.pmem[7587] ;
wire \u_lsu.pmem[7588] ;
wire \u_lsu.pmem[7589] ;
wire \u_lsu.pmem[7590] ;
wire \u_lsu.pmem[7591] ;
wire \u_lsu.pmem[7592] ;
wire \u_lsu.pmem[7593] ;
wire \u_lsu.pmem[7594] ;
wire \u_lsu.pmem[7595] ;
wire \u_lsu.pmem[7596] ;
wire \u_lsu.pmem[7597] ;
wire \u_lsu.pmem[7598] ;
wire \u_lsu.pmem[7599] ;
wire \u_lsu.pmem[7600] ;
wire \u_lsu.pmem[7601] ;
wire \u_lsu.pmem[7602] ;
wire \u_lsu.pmem[7603] ;
wire \u_lsu.pmem[7604] ;
wire \u_lsu.pmem[7605] ;
wire \u_lsu.pmem[7606] ;
wire \u_lsu.pmem[7607] ;
wire \u_lsu.pmem[7608] ;
wire \u_lsu.pmem[7609] ;
wire \u_lsu.pmem[7610] ;
wire \u_lsu.pmem[7611] ;
wire \u_lsu.pmem[7612] ;
wire \u_lsu.pmem[7613] ;
wire \u_lsu.pmem[7614] ;
wire \u_lsu.pmem[7615] ;
wire \u_lsu.pmem[7616] ;
wire \u_lsu.pmem[7617] ;
wire \u_lsu.pmem[7618] ;
wire \u_lsu.pmem[7619] ;
wire \u_lsu.pmem[7620] ;
wire \u_lsu.pmem[7621] ;
wire \u_lsu.pmem[7622] ;
wire \u_lsu.pmem[7623] ;
wire \u_lsu.pmem[7624] ;
wire \u_lsu.pmem[7625] ;
wire \u_lsu.pmem[7626] ;
wire \u_lsu.pmem[7627] ;
wire \u_lsu.pmem[7628] ;
wire \u_lsu.pmem[7629] ;
wire \u_lsu.pmem[7630] ;
wire \u_lsu.pmem[7631] ;
wire \u_lsu.pmem[7632] ;
wire \u_lsu.pmem[7633] ;
wire \u_lsu.pmem[7634] ;
wire \u_lsu.pmem[7635] ;
wire \u_lsu.pmem[7636] ;
wire \u_lsu.pmem[7637] ;
wire \u_lsu.pmem[7638] ;
wire \u_lsu.pmem[7639] ;
wire \u_lsu.pmem[7640] ;
wire \u_lsu.pmem[7641] ;
wire \u_lsu.pmem[7642] ;
wire \u_lsu.pmem[7643] ;
wire \u_lsu.pmem[7644] ;
wire \u_lsu.pmem[7645] ;
wire \u_lsu.pmem[7646] ;
wire \u_lsu.pmem[7647] ;
wire \u_lsu.pmem[7648] ;
wire \u_lsu.pmem[7649] ;
wire \u_lsu.pmem[7650] ;
wire \u_lsu.pmem[7651] ;
wire \u_lsu.pmem[7652] ;
wire \u_lsu.pmem[7653] ;
wire \u_lsu.pmem[7654] ;
wire \u_lsu.pmem[7655] ;
wire \u_lsu.pmem[7656] ;
wire \u_lsu.pmem[7657] ;
wire \u_lsu.pmem[7658] ;
wire \u_lsu.pmem[7659] ;
wire \u_lsu.pmem[7660] ;
wire \u_lsu.pmem[7661] ;
wire \u_lsu.pmem[7662] ;
wire \u_lsu.pmem[7663] ;
wire \u_lsu.pmem[7664] ;
wire \u_lsu.pmem[7665] ;
wire \u_lsu.pmem[7666] ;
wire \u_lsu.pmem[7667] ;
wire \u_lsu.pmem[7668] ;
wire \u_lsu.pmem[7669] ;
wire \u_lsu.pmem[7670] ;
wire \u_lsu.pmem[7671] ;
wire \u_lsu.pmem[7672] ;
wire \u_lsu.pmem[7673] ;
wire \u_lsu.pmem[7674] ;
wire \u_lsu.pmem[7675] ;
wire \u_lsu.pmem[7676] ;
wire \u_lsu.pmem[7677] ;
wire \u_lsu.pmem[7678] ;
wire \u_lsu.pmem[7679] ;
wire \u_lsu.pmem[7680] ;
wire \u_lsu.pmem[7681] ;
wire \u_lsu.pmem[7682] ;
wire \u_lsu.pmem[7683] ;
wire \u_lsu.pmem[7684] ;
wire \u_lsu.pmem[7685] ;
wire \u_lsu.pmem[7686] ;
wire \u_lsu.pmem[7687] ;
wire \u_lsu.pmem[7688] ;
wire \u_lsu.pmem[7689] ;
wire \u_lsu.pmem[7690] ;
wire \u_lsu.pmem[7691] ;
wire \u_lsu.pmem[7692] ;
wire \u_lsu.pmem[7693] ;
wire \u_lsu.pmem[7694] ;
wire \u_lsu.pmem[7695] ;
wire \u_lsu.pmem[7696] ;
wire \u_lsu.pmem[7697] ;
wire \u_lsu.pmem[7698] ;
wire \u_lsu.pmem[7699] ;
wire \u_lsu.pmem[7700] ;
wire \u_lsu.pmem[7701] ;
wire \u_lsu.pmem[7702] ;
wire \u_lsu.pmem[7703] ;
wire \u_lsu.pmem[7704] ;
wire \u_lsu.pmem[7705] ;
wire \u_lsu.pmem[7706] ;
wire \u_lsu.pmem[7707] ;
wire \u_lsu.pmem[7708] ;
wire \u_lsu.pmem[7709] ;
wire \u_lsu.pmem[7710] ;
wire \u_lsu.pmem[7711] ;
wire \u_lsu.pmem[7712] ;
wire \u_lsu.pmem[7713] ;
wire \u_lsu.pmem[7714] ;
wire \u_lsu.pmem[7715] ;
wire \u_lsu.pmem[7716] ;
wire \u_lsu.pmem[7717] ;
wire \u_lsu.pmem[7718] ;
wire \u_lsu.pmem[7719] ;
wire \u_lsu.pmem[7720] ;
wire \u_lsu.pmem[7721] ;
wire \u_lsu.pmem[7722] ;
wire \u_lsu.pmem[7723] ;
wire \u_lsu.pmem[7724] ;
wire \u_lsu.pmem[7725] ;
wire \u_lsu.pmem[7726] ;
wire \u_lsu.pmem[7727] ;
wire \u_lsu.pmem[7728] ;
wire \u_lsu.pmem[7729] ;
wire \u_lsu.pmem[7730] ;
wire \u_lsu.pmem[7731] ;
wire \u_lsu.pmem[7732] ;
wire \u_lsu.pmem[7733] ;
wire \u_lsu.pmem[7734] ;
wire \u_lsu.pmem[7735] ;
wire \u_lsu.pmem[7736] ;
wire \u_lsu.pmem[7737] ;
wire \u_lsu.pmem[7738] ;
wire \u_lsu.pmem[7739] ;
wire \u_lsu.pmem[7740] ;
wire \u_lsu.pmem[7741] ;
wire \u_lsu.pmem[7742] ;
wire \u_lsu.pmem[7743] ;
wire \u_lsu.pmem[7744] ;
wire \u_lsu.pmem[7745] ;
wire \u_lsu.pmem[7746] ;
wire \u_lsu.pmem[7747] ;
wire \u_lsu.pmem[7748] ;
wire \u_lsu.pmem[7749] ;
wire \u_lsu.pmem[7750] ;
wire \u_lsu.pmem[7751] ;
wire \u_lsu.pmem[7752] ;
wire \u_lsu.pmem[7753] ;
wire \u_lsu.pmem[7754] ;
wire \u_lsu.pmem[7755] ;
wire \u_lsu.pmem[7756] ;
wire \u_lsu.pmem[7757] ;
wire \u_lsu.pmem[7758] ;
wire \u_lsu.pmem[7759] ;
wire \u_lsu.pmem[7760] ;
wire \u_lsu.pmem[7761] ;
wire \u_lsu.pmem[7762] ;
wire \u_lsu.pmem[7763] ;
wire \u_lsu.pmem[7764] ;
wire \u_lsu.pmem[7765] ;
wire \u_lsu.pmem[7766] ;
wire \u_lsu.pmem[7767] ;
wire \u_lsu.pmem[7768] ;
wire \u_lsu.pmem[7769] ;
wire \u_lsu.pmem[7770] ;
wire \u_lsu.pmem[7771] ;
wire \u_lsu.pmem[7772] ;
wire \u_lsu.pmem[7773] ;
wire \u_lsu.pmem[7774] ;
wire \u_lsu.pmem[7775] ;
wire \u_lsu.pmem[7776] ;
wire \u_lsu.pmem[7777] ;
wire \u_lsu.pmem[7778] ;
wire \u_lsu.pmem[7779] ;
wire \u_lsu.pmem[7780] ;
wire \u_lsu.pmem[7781] ;
wire \u_lsu.pmem[7782] ;
wire \u_lsu.pmem[7783] ;
wire \u_lsu.pmem[7784] ;
wire \u_lsu.pmem[7785] ;
wire \u_lsu.pmem[7786] ;
wire \u_lsu.pmem[7787] ;
wire \u_lsu.pmem[7788] ;
wire \u_lsu.pmem[7789] ;
wire \u_lsu.pmem[7790] ;
wire \u_lsu.pmem[7791] ;
wire \u_lsu.pmem[7792] ;
wire \u_lsu.pmem[7793] ;
wire \u_lsu.pmem[7794] ;
wire \u_lsu.pmem[7795] ;
wire \u_lsu.pmem[7796] ;
wire \u_lsu.pmem[7797] ;
wire \u_lsu.pmem[7798] ;
wire \u_lsu.pmem[7799] ;
wire \u_lsu.pmem[7800] ;
wire \u_lsu.pmem[7801] ;
wire \u_lsu.pmem[7802] ;
wire \u_lsu.pmem[7803] ;
wire \u_lsu.pmem[7804] ;
wire \u_lsu.pmem[7805] ;
wire \u_lsu.pmem[7806] ;
wire \u_lsu.pmem[7807] ;
wire \u_lsu.pmem[7808] ;
wire \u_lsu.pmem[7809] ;
wire \u_lsu.pmem[7810] ;
wire \u_lsu.pmem[7811] ;
wire \u_lsu.pmem[7812] ;
wire \u_lsu.pmem[7813] ;
wire \u_lsu.pmem[7814] ;
wire \u_lsu.pmem[7815] ;
wire \u_lsu.pmem[7816] ;
wire \u_lsu.pmem[7817] ;
wire \u_lsu.pmem[7818] ;
wire \u_lsu.pmem[7819] ;
wire \u_lsu.pmem[7820] ;
wire \u_lsu.pmem[7821] ;
wire \u_lsu.pmem[7822] ;
wire \u_lsu.pmem[7823] ;
wire \u_lsu.pmem[7824] ;
wire \u_lsu.pmem[7825] ;
wire \u_lsu.pmem[7826] ;
wire \u_lsu.pmem[7827] ;
wire \u_lsu.pmem[7828] ;
wire \u_lsu.pmem[7829] ;
wire \u_lsu.pmem[7830] ;
wire \u_lsu.pmem[7831] ;
wire \u_lsu.pmem[7832] ;
wire \u_lsu.pmem[7833] ;
wire \u_lsu.pmem[7834] ;
wire \u_lsu.pmem[7835] ;
wire \u_lsu.pmem[7836] ;
wire \u_lsu.pmem[7837] ;
wire \u_lsu.pmem[7838] ;
wire \u_lsu.pmem[7839] ;
wire \u_lsu.pmem[7840] ;
wire \u_lsu.pmem[7841] ;
wire \u_lsu.pmem[7842] ;
wire \u_lsu.pmem[7843] ;
wire \u_lsu.pmem[7844] ;
wire \u_lsu.pmem[7845] ;
wire \u_lsu.pmem[7846] ;
wire \u_lsu.pmem[7847] ;
wire \u_lsu.pmem[7848] ;
wire \u_lsu.pmem[7849] ;
wire \u_lsu.pmem[7850] ;
wire \u_lsu.pmem[7851] ;
wire \u_lsu.pmem[7852] ;
wire \u_lsu.pmem[7853] ;
wire \u_lsu.pmem[7854] ;
wire \u_lsu.pmem[7855] ;
wire \u_lsu.pmem[7856] ;
wire \u_lsu.pmem[7857] ;
wire \u_lsu.pmem[7858] ;
wire \u_lsu.pmem[7859] ;
wire \u_lsu.pmem[7860] ;
wire \u_lsu.pmem[7861] ;
wire \u_lsu.pmem[7862] ;
wire \u_lsu.pmem[7863] ;
wire \u_lsu.pmem[7864] ;
wire \u_lsu.pmem[7865] ;
wire \u_lsu.pmem[7866] ;
wire \u_lsu.pmem[7867] ;
wire \u_lsu.pmem[7868] ;
wire \u_lsu.pmem[7869] ;
wire \u_lsu.pmem[7870] ;
wire \u_lsu.pmem[7871] ;
wire \u_lsu.pmem[7872] ;
wire \u_lsu.pmem[7873] ;
wire \u_lsu.pmem[7874] ;
wire \u_lsu.pmem[7875] ;
wire \u_lsu.pmem[7876] ;
wire \u_lsu.pmem[7877] ;
wire \u_lsu.pmem[7878] ;
wire \u_lsu.pmem[7879] ;
wire \u_lsu.pmem[7880] ;
wire \u_lsu.pmem[7881] ;
wire \u_lsu.pmem[7882] ;
wire \u_lsu.pmem[7883] ;
wire \u_lsu.pmem[7884] ;
wire \u_lsu.pmem[7885] ;
wire \u_lsu.pmem[7886] ;
wire \u_lsu.pmem[7887] ;
wire \u_lsu.pmem[7888] ;
wire \u_lsu.pmem[7889] ;
wire \u_lsu.pmem[7890] ;
wire \u_lsu.pmem[7891] ;
wire \u_lsu.pmem[7892] ;
wire \u_lsu.pmem[7893] ;
wire \u_lsu.pmem[7894] ;
wire \u_lsu.pmem[7895] ;
wire \u_lsu.pmem[7896] ;
wire \u_lsu.pmem[7897] ;
wire \u_lsu.pmem[7898] ;
wire \u_lsu.pmem[7899] ;
wire \u_lsu.pmem[7900] ;
wire \u_lsu.pmem[7901] ;
wire \u_lsu.pmem[7902] ;
wire \u_lsu.pmem[7903] ;
wire \u_lsu.pmem[7904] ;
wire \u_lsu.pmem[7905] ;
wire \u_lsu.pmem[7906] ;
wire \u_lsu.pmem[7907] ;
wire \u_lsu.pmem[7908] ;
wire \u_lsu.pmem[7909] ;
wire \u_lsu.pmem[7910] ;
wire \u_lsu.pmem[7911] ;
wire \u_lsu.pmem[7912] ;
wire \u_lsu.pmem[7913] ;
wire \u_lsu.pmem[7914] ;
wire \u_lsu.pmem[7915] ;
wire \u_lsu.pmem[7916] ;
wire \u_lsu.pmem[7917] ;
wire \u_lsu.pmem[7918] ;
wire \u_lsu.pmem[7919] ;
wire \u_lsu.pmem[7920] ;
wire \u_lsu.pmem[7921] ;
wire \u_lsu.pmem[7922] ;
wire \u_lsu.pmem[7923] ;
wire \u_lsu.pmem[7924] ;
wire \u_lsu.pmem[7925] ;
wire \u_lsu.pmem[7926] ;
wire \u_lsu.pmem[7927] ;
wire \u_lsu.pmem[7928] ;
wire \u_lsu.pmem[7929] ;
wire \u_lsu.pmem[7930] ;
wire \u_lsu.pmem[7931] ;
wire \u_lsu.pmem[7932] ;
wire \u_lsu.pmem[7933] ;
wire \u_lsu.pmem[7934] ;
wire \u_lsu.pmem[7935] ;
wire \u_lsu.pmem[7936] ;
wire \u_lsu.pmem[7937] ;
wire \u_lsu.pmem[7938] ;
wire \u_lsu.pmem[7939] ;
wire \u_lsu.pmem[7940] ;
wire \u_lsu.pmem[7941] ;
wire \u_lsu.pmem[7942] ;
wire \u_lsu.pmem[7943] ;
wire \u_lsu.pmem[7944] ;
wire \u_lsu.pmem[7945] ;
wire \u_lsu.pmem[7946] ;
wire \u_lsu.pmem[7947] ;
wire \u_lsu.pmem[7948] ;
wire \u_lsu.pmem[7949] ;
wire \u_lsu.pmem[7950] ;
wire \u_lsu.pmem[7951] ;
wire \u_lsu.pmem[7952] ;
wire \u_lsu.pmem[7953] ;
wire \u_lsu.pmem[7954] ;
wire \u_lsu.pmem[7955] ;
wire \u_lsu.pmem[7956] ;
wire \u_lsu.pmem[7957] ;
wire \u_lsu.pmem[7958] ;
wire \u_lsu.pmem[7959] ;
wire \u_lsu.pmem[7960] ;
wire \u_lsu.pmem[7961] ;
wire \u_lsu.pmem[7962] ;
wire \u_lsu.pmem[7963] ;
wire \u_lsu.pmem[7964] ;
wire \u_lsu.pmem[7965] ;
wire \u_lsu.pmem[7966] ;
wire \u_lsu.pmem[7967] ;
wire \u_lsu.pmem[7968] ;
wire \u_lsu.pmem[7969] ;
wire \u_lsu.pmem[7970] ;
wire \u_lsu.pmem[7971] ;
wire \u_lsu.pmem[7972] ;
wire \u_lsu.pmem[7973] ;
wire \u_lsu.pmem[7974] ;
wire \u_lsu.pmem[7975] ;
wire \u_lsu.pmem[7976] ;
wire \u_lsu.pmem[7977] ;
wire \u_lsu.pmem[7978] ;
wire \u_lsu.pmem[7979] ;
wire \u_lsu.pmem[7980] ;
wire \u_lsu.pmem[7981] ;
wire \u_lsu.pmem[7982] ;
wire \u_lsu.pmem[7983] ;
wire \u_lsu.pmem[7984] ;
wire \u_lsu.pmem[7985] ;
wire \u_lsu.pmem[7986] ;
wire \u_lsu.pmem[7987] ;
wire \u_lsu.pmem[7988] ;
wire \u_lsu.pmem[7989] ;
wire \u_lsu.pmem[7990] ;
wire \u_lsu.pmem[7991] ;
wire \u_lsu.pmem[7992] ;
wire \u_lsu.pmem[7993] ;
wire \u_lsu.pmem[7994] ;
wire \u_lsu.pmem[7995] ;
wire \u_lsu.pmem[7996] ;
wire \u_lsu.pmem[7997] ;
wire \u_lsu.pmem[7998] ;
wire \u_lsu.pmem[7999] ;
wire \u_lsu.pmem[8000] ;
wire \u_lsu.pmem[8001] ;
wire \u_lsu.pmem[8002] ;
wire \u_lsu.pmem[8003] ;
wire \u_lsu.pmem[8004] ;
wire \u_lsu.pmem[8005] ;
wire \u_lsu.pmem[8006] ;
wire \u_lsu.pmem[8007] ;
wire \u_lsu.pmem[8008] ;
wire \u_lsu.pmem[8009] ;
wire \u_lsu.pmem[8010] ;
wire \u_lsu.pmem[8011] ;
wire \u_lsu.pmem[8012] ;
wire \u_lsu.pmem[8013] ;
wire \u_lsu.pmem[8014] ;
wire \u_lsu.pmem[8015] ;
wire \u_lsu.pmem[8016] ;
wire \u_lsu.pmem[8017] ;
wire \u_lsu.pmem[8018] ;
wire \u_lsu.pmem[8019] ;
wire \u_lsu.pmem[8020] ;
wire \u_lsu.pmem[8021] ;
wire \u_lsu.pmem[8022] ;
wire \u_lsu.pmem[8023] ;
wire \u_lsu.pmem[8024] ;
wire \u_lsu.pmem[8025] ;
wire \u_lsu.pmem[8026] ;
wire \u_lsu.pmem[8027] ;
wire \u_lsu.pmem[8028] ;
wire \u_lsu.pmem[8029] ;
wire \u_lsu.pmem[8030] ;
wire \u_lsu.pmem[8031] ;
wire \u_lsu.pmem[8032] ;
wire \u_lsu.pmem[8033] ;
wire \u_lsu.pmem[8034] ;
wire \u_lsu.pmem[8035] ;
wire \u_lsu.pmem[8036] ;
wire \u_lsu.pmem[8037] ;
wire \u_lsu.pmem[8038] ;
wire \u_lsu.pmem[8039] ;
wire \u_lsu.pmem[8040] ;
wire \u_lsu.pmem[8041] ;
wire \u_lsu.pmem[8042] ;
wire \u_lsu.pmem[8043] ;
wire \u_lsu.pmem[8044] ;
wire \u_lsu.pmem[8045] ;
wire \u_lsu.pmem[8046] ;
wire \u_lsu.pmem[8047] ;
wire \u_lsu.pmem[8048] ;
wire \u_lsu.pmem[8049] ;
wire \u_lsu.pmem[8050] ;
wire \u_lsu.pmem[8051] ;
wire \u_lsu.pmem[8052] ;
wire \u_lsu.pmem[8053] ;
wire \u_lsu.pmem[8054] ;
wire \u_lsu.pmem[8055] ;
wire \u_lsu.pmem[8056] ;
wire \u_lsu.pmem[8057] ;
wire \u_lsu.pmem[8058] ;
wire \u_lsu.pmem[8059] ;
wire \u_lsu.pmem[8060] ;
wire \u_lsu.pmem[8061] ;
wire \u_lsu.pmem[8062] ;
wire \u_lsu.pmem[8063] ;
wire \u_lsu.pmem[8064] ;
wire \u_lsu.pmem[8065] ;
wire \u_lsu.pmem[8066] ;
wire \u_lsu.pmem[8067] ;
wire \u_lsu.pmem[8068] ;
wire \u_lsu.pmem[8069] ;
wire \u_lsu.pmem[8070] ;
wire \u_lsu.pmem[8071] ;
wire \u_lsu.pmem[8072] ;
wire \u_lsu.pmem[8073] ;
wire \u_lsu.pmem[8074] ;
wire \u_lsu.pmem[8075] ;
wire \u_lsu.pmem[8076] ;
wire \u_lsu.pmem[8077] ;
wire \u_lsu.pmem[8078] ;
wire \u_lsu.pmem[8079] ;
wire \u_lsu.pmem[8080] ;
wire \u_lsu.pmem[8081] ;
wire \u_lsu.pmem[8082] ;
wire \u_lsu.pmem[8083] ;
wire \u_lsu.pmem[8084] ;
wire \u_lsu.pmem[8085] ;
wire \u_lsu.pmem[8086] ;
wire \u_lsu.pmem[8087] ;
wire \u_lsu.pmem[8088] ;
wire \u_lsu.pmem[8089] ;
wire \u_lsu.pmem[8090] ;
wire \u_lsu.pmem[8091] ;
wire \u_lsu.pmem[8092] ;
wire \u_lsu.pmem[8093] ;
wire \u_lsu.pmem[8094] ;
wire \u_lsu.pmem[8095] ;
wire \u_lsu.pmem[8096] ;
wire \u_lsu.pmem[8097] ;
wire \u_lsu.pmem[8098] ;
wire \u_lsu.pmem[8099] ;
wire \u_lsu.pmem[8100] ;
wire \u_lsu.pmem[8101] ;
wire \u_lsu.pmem[8102] ;
wire \u_lsu.pmem[8103] ;
wire \u_lsu.pmem[8104] ;
wire \u_lsu.pmem[8105] ;
wire \u_lsu.pmem[8106] ;
wire \u_lsu.pmem[8107] ;
wire \u_lsu.pmem[8108] ;
wire \u_lsu.pmem[8109] ;
wire \u_lsu.pmem[8110] ;
wire \u_lsu.pmem[8111] ;
wire \u_lsu.pmem[8112] ;
wire \u_lsu.pmem[8113] ;
wire \u_lsu.pmem[8114] ;
wire \u_lsu.pmem[8115] ;
wire \u_lsu.pmem[8116] ;
wire \u_lsu.pmem[8117] ;
wire \u_lsu.pmem[8118] ;
wire \u_lsu.pmem[8119] ;
wire \u_lsu.pmem[8120] ;
wire \u_lsu.pmem[8121] ;
wire \u_lsu.pmem[8122] ;
wire \u_lsu.pmem[8123] ;
wire \u_lsu.pmem[8124] ;
wire \u_lsu.pmem[8125] ;
wire \u_lsu.pmem[8126] ;
wire \u_lsu.pmem[8127] ;
wire \u_lsu.pmem[8128] ;
wire \u_lsu.pmem[8129] ;
wire \u_lsu.pmem[8130] ;
wire \u_lsu.pmem[8131] ;
wire \u_lsu.pmem[8132] ;
wire \u_lsu.pmem[8133] ;
wire \u_lsu.pmem[8134] ;
wire \u_lsu.pmem[8135] ;
wire \u_lsu.pmem[8136] ;
wire \u_lsu.pmem[8137] ;
wire \u_lsu.pmem[8138] ;
wire \u_lsu.pmem[8139] ;
wire \u_lsu.pmem[8140] ;
wire \u_lsu.pmem[8141] ;
wire \u_lsu.pmem[8142] ;
wire \u_lsu.pmem[8143] ;
wire \u_lsu.pmem[8144] ;
wire \u_lsu.pmem[8145] ;
wire \u_lsu.pmem[8146] ;
wire \u_lsu.pmem[8147] ;
wire \u_lsu.pmem[8148] ;
wire \u_lsu.pmem[8149] ;
wire \u_lsu.pmem[8150] ;
wire \u_lsu.pmem[8151] ;
wire \u_lsu.pmem[8152] ;
wire \u_lsu.pmem[8153] ;
wire \u_lsu.pmem[8154] ;
wire \u_lsu.pmem[8155] ;
wire \u_lsu.pmem[8156] ;
wire \u_lsu.pmem[8157] ;
wire \u_lsu.pmem[8158] ;
wire \u_lsu.pmem[8159] ;
wire \u_lsu.pmem[8160] ;
wire \u_lsu.pmem[8161] ;
wire \u_lsu.pmem[8162] ;
wire \u_lsu.pmem[8163] ;
wire \u_lsu.pmem[8164] ;
wire \u_lsu.pmem[8165] ;
wire \u_lsu.pmem[8166] ;
wire \u_lsu.pmem[8167] ;

assign alu_result_out[0] = \alu_result_out[0] ;
assign alu_result_out[1] = \alu_result_out[1] ;
assign alu_result_out[2] = \alu_result_out[2] ;
assign alu_result_out[3] = \alu_result_out[3] ;
assign alu_result_out[4] = \alu_result_out[4] ;
assign alu_result_out[5] = \alu_result_out[5] ;
assign alu_result_out[6] = \alu_result_out[6] ;
assign alu_result_out[7] = \alu_result_out[7] ;
assign alu_result_out[8] = \alu_result_out[8] ;
assign alu_result_out[9] = \alu_result_out[9] ;
assign alu_result_out[10] = \alu_result_out[10] ;
assign alu_result_out[11] = \alu_result_out[11] ;
assign alu_result_out[12] = \alu_result_out[12] ;
assign alu_result_out[13] = \alu_result_out[13] ;
assign alu_result_out[14] = \alu_result_out[14] ;
assign alu_result_out[15] = \alu_result_out[15] ;
assign alu_result_out[16] = \alu_result_out[16] ;
assign alu_result_out[17] = \alu_result_out[17] ;
assign alu_result_out[18] = \alu_result_out[18] ;
assign alu_result_out[19] = \alu_result_out[19] ;
assign alu_result_out[20] = \alu_result_out[20] ;
assign alu_result_out[21] = \alu_result_out[21] ;
assign alu_result_out[22] = \alu_result_out[22] ;
assign alu_result_out[23] = \alu_result_out[23] ;
assign alu_result_out[24] = \alu_result_out[24] ;
assign alu_result_out[25] = \alu_result_out[25] ;
assign alu_result_out[26] = \alu_result_out[26] ;
assign alu_result_out[27] = \alu_result_out[27] ;
assign alu_result_out[28] = \alu_result_out[28] ;
assign alu_result_out[29] = \alu_result_out[29] ;
assign alu_result_out[30] = \alu_result_out[30] ;
assign alu_result_out[31] = \alu_result_out[31] ;
assign load_data_out[0] = \load_data_out[0] ;
assign load_data_out[1] = \load_data_out[1] ;
assign load_data_out[2] = \load_data_out[2] ;
assign load_data_out[3] = \load_data_out[3] ;
assign load_data_out[4] = \load_data_out[4] ;
assign load_data_out[5] = \load_data_out[5] ;
assign load_data_out[6] = \load_data_out[6] ;
assign load_data_out[10] = \load_data_out[7] ;
assign load_data_out[10] = \load_data_out[8] ;
assign load_data_out[10] = \load_data_out[9] ;
assign load_data_out[10] = \load_data_out[10] ;
assign load_data_out[10] = \load_data_out[11] ;
assign load_data_out[10] = \load_data_out[12] ;
assign load_data_out[10] = \load_data_out[13] ;
assign load_data_out[10] = \load_data_out[14] ;
assign load_data_out[10] = \load_data_out[15] ;
assign load_data_out[10] = \load_data_out[16] ;
assign load_data_out[10] = \load_data_out[17] ;
assign load_data_out[10] = \load_data_out[18] ;
assign load_data_out[10] = \load_data_out[19] ;
assign load_data_out[10] = \load_data_out[20] ;
assign load_data_out[10] = \load_data_out[21] ;
assign load_data_out[10] = \load_data_out[22] ;
assign load_data_out[10] = \load_data_out[23] ;
assign load_data_out[10] = \load_data_out[24] ;
assign load_data_out[10] = \load_data_out[25] ;
assign load_data_out[10] = \load_data_out[26] ;
assign load_data_out[10] = \load_data_out[27] ;
assign load_data_out[10] = \load_data_out[28] ;
assign load_data_out[10] = \load_data_out[29] ;
assign load_data_out[10] = \load_data_out[30] ;
assign load_data_out[10] = \load_data_out[31] ;
assign pc_out[0] = \pc_out[0] ;
assign pc_out[1] = \pc_out[1] ;
assign pc_out[2] = \pc_out[2] ;
assign pc_out[3] = \pc_out[3] ;
assign pc_out[4] = \pc_out[4] ;
assign pc_out[5] = \pc_out[5] ;
assign pc_out[6] = \pc_out[6] ;
assign pc_out[7] = \pc_out[7] ;
assign pc_out[8] = \pc_out[8] ;
assign pc_out[9] = \pc_out[9] ;
assign pc_out[10] = \pc_out[10] ;
assign pc_out[11] = \pc_out[11] ;
assign pc_out[12] = \pc_out[12] ;
assign pc_out[13] = \pc_out[13] ;
assign pc_out[14] = \pc_out[14] ;
assign pc_out[15] = \pc_out[15] ;
assign pc_out[16] = \pc_out[16] ;
assign pc_out[17] = \pc_out[17] ;
assign pc_out[18] = \pc_out[18] ;
assign pc_out[19] = \pc_out[19] ;
assign pc_out[20] = \pc_out[20] ;
assign pc_out[21] = \pc_out[21] ;
assign pc_out[22] = \pc_out[22] ;
assign pc_out[23] = \pc_out[23] ;
assign pc_out[24] = \pc_out[24] ;
assign pc_out[25] = \pc_out[25] ;
assign pc_out[26] = \pc_out[26] ;
assign pc_out[27] = \pc_out[27] ;
assign pc_out[28] = \pc_out[28] ;
assign pc_out[29] = \pc_out[29] ;
assign pc_out[30] = \pc_out[30] ;
assign pc_out[31] = \pc_out[31] ;

INV_X1 _12022_ ( .A(dnpc_$_NOT__Y_A_$_ANDNOT__B_A ), .ZN(_08575_ ) );
MUX2_X1 _12023_ ( .A(\u_gpr.regfile[0][7] ), .B(\u_gpr.regfile[1][7] ), .S(fanout_net_5 ), .Z(_08576_ ) );
MUX2_X1 _12024_ ( .A(\u_gpr.regfile[2][7] ), .B(\u_gpr.regfile[3][7] ), .S(fanout_net_5 ), .Z(_08577_ ) );
MUX2_X1 _12025_ ( .A(_08576_ ), .B(_08577_ ), .S(fanout_net_7 ), .Z(_08578_ ) );
NOR2_X1 _12026_ ( .A1(fanout_net_7 ), .A2(fanout_net_5 ), .ZN(_08579_ ) );
INV_X1 _12027_ ( .A(_08579_ ), .ZN(_08580_ ) );
AND2_X1 _12028_ ( .A1(_08578_ ), .A2(_08580_ ), .ZN(_08581_ ) );
BUF_X4 _12029_ ( .A(_08581_ ), .Z(_08582_ ) );
MUX2_X1 _12030_ ( .A(\u_gpr.regfile[0][7] ), .B(\u_gpr.regfile[1][7] ), .S(fanout_net_2 ), .Z(_08583_ ) );
MUX2_X1 _12031_ ( .A(\u_gpr.regfile[2][7] ), .B(\u_gpr.regfile[3][7] ), .S(fanout_net_2 ), .Z(_08584_ ) );
MUX2_X1 _12032_ ( .A(_08583_ ), .B(_08584_ ), .S(fanout_net_4 ), .Z(_08585_ ) );
INV_X1 _12033_ ( .A(fanout_net_4 ), .ZN(_08586_ ) );
INV_X1 _12034_ ( .A(fanout_net_2 ), .ZN(_08587_ ) );
NAND2_X1 _12035_ ( .A1(_08586_ ), .A2(_08587_ ), .ZN(_08588_ ) );
CLKBUF_X2 _12036_ ( .A(_08588_ ), .Z(_08589_ ) );
AND2_X1 _12037_ ( .A1(_08585_ ), .A2(_08589_ ), .ZN(_08590_ ) );
XNOR2_X1 _12038_ ( .A(_08582_ ), .B(_08590_ ), .ZN(_08591_ ) );
MUX2_X1 _12039_ ( .A(\u_gpr.regfile[0][5] ), .B(\u_gpr.regfile[1][5] ), .S(fanout_net_5 ), .Z(_08592_ ) );
MUX2_X1 _12040_ ( .A(\u_gpr.regfile[2][5] ), .B(\u_gpr.regfile[3][5] ), .S(fanout_net_5 ), .Z(_08593_ ) );
MUX2_X1 _12041_ ( .A(_08592_ ), .B(_08593_ ), .S(fanout_net_7 ), .Z(_08594_ ) );
AND2_X1 _12042_ ( .A1(_08594_ ), .A2(_08580_ ), .ZN(_08595_ ) );
MUX2_X1 _12043_ ( .A(\u_gpr.regfile[0][5] ), .B(\u_gpr.regfile[1][5] ), .S(fanout_net_2 ), .Z(_08596_ ) );
MUX2_X1 _12044_ ( .A(\u_gpr.regfile[2][5] ), .B(\u_gpr.regfile[3][5] ), .S(fanout_net_2 ), .Z(_08597_ ) );
MUX2_X1 _12045_ ( .A(_08596_ ), .B(_08597_ ), .S(fanout_net_4 ), .Z(_08598_ ) );
AND2_X1 _12046_ ( .A1(_08598_ ), .A2(_08589_ ), .ZN(_08599_ ) );
XNOR2_X1 _12047_ ( .A(_08595_ ), .B(_08599_ ), .ZN(_08600_ ) );
MUX2_X1 _12048_ ( .A(\u_gpr.regfile[0][4] ), .B(\u_gpr.regfile[1][4] ), .S(fanout_net_5 ), .Z(_08601_ ) );
MUX2_X1 _12049_ ( .A(\u_gpr.regfile[2][4] ), .B(\u_gpr.regfile[3][4] ), .S(fanout_net_5 ), .Z(_08602_ ) );
MUX2_X1 _12050_ ( .A(_08601_ ), .B(_08602_ ), .S(fanout_net_7 ), .Z(_08603_ ) );
AND2_X1 _12051_ ( .A1(_08603_ ), .A2(_08580_ ), .ZN(_08604_ ) );
BUF_X4 _12052_ ( .A(_08604_ ), .Z(_08605_ ) );
MUX2_X1 _12053_ ( .A(\u_gpr.regfile[0][4] ), .B(\u_gpr.regfile[1][4] ), .S(fanout_net_2 ), .Z(_08606_ ) );
MUX2_X1 _12054_ ( .A(\u_gpr.regfile[2][4] ), .B(\u_gpr.regfile[3][4] ), .S(fanout_net_2 ), .Z(_08607_ ) );
MUX2_X1 _12055_ ( .A(_08606_ ), .B(_08607_ ), .S(fanout_net_4 ), .Z(_08608_ ) );
CLKBUF_X2 _12056_ ( .A(_08589_ ), .Z(_08609_ ) );
CLKBUF_X2 _12057_ ( .A(_08609_ ), .Z(_08610_ ) );
BUF_X2 _12058_ ( .A(_08610_ ), .Z(_08611_ ) );
AND2_X1 _12059_ ( .A1(_08608_ ), .A2(_08611_ ), .ZN(_08612_ ) );
XNOR2_X1 _12060_ ( .A(_08605_ ), .B(_08612_ ), .ZN(_08613_ ) );
MUX2_X1 _12061_ ( .A(\u_gpr.regfile[0][6] ), .B(\u_gpr.regfile[1][6] ), .S(fanout_net_5 ), .Z(_08614_ ) );
MUX2_X1 _12062_ ( .A(\u_gpr.regfile[2][6] ), .B(\u_gpr.regfile[3][6] ), .S(fanout_net_5 ), .Z(_08615_ ) );
MUX2_X1 _12063_ ( .A(_08614_ ), .B(_08615_ ), .S(fanout_net_7 ), .Z(_08616_ ) );
AND2_X1 _12064_ ( .A1(_08616_ ), .A2(_08580_ ), .ZN(_08617_ ) );
MUX2_X1 _12065_ ( .A(\u_gpr.regfile[0][6] ), .B(\u_gpr.regfile[1][6] ), .S(fanout_net_2 ), .Z(_08618_ ) );
MUX2_X1 _12066_ ( .A(\u_gpr.regfile[2][6] ), .B(\u_gpr.regfile[3][6] ), .S(fanout_net_2 ), .Z(_08619_ ) );
MUX2_X1 _12067_ ( .A(_08618_ ), .B(_08619_ ), .S(fanout_net_4 ), .Z(_08620_ ) );
AND2_X1 _12068_ ( .A1(_08620_ ), .A2(_08589_ ), .ZN(_08621_ ) );
XNOR2_X1 _12069_ ( .A(_08617_ ), .B(_08621_ ), .ZN(_08622_ ) );
NAND4_X1 _12070_ ( .A1(_08591_ ), .A2(_08600_ ), .A3(_08613_ ), .A4(_08622_ ), .ZN(_08623_ ) );
MUX2_X1 _12071_ ( .A(\u_gpr.regfile[0][0] ), .B(\u_gpr.regfile[1][0] ), .S(fanout_net_2 ), .Z(_08624_ ) );
MUX2_X1 _12072_ ( .A(\u_gpr.regfile[2][0] ), .B(\u_gpr.regfile[3][0] ), .S(fanout_net_2 ), .Z(_08625_ ) );
MUX2_X1 _12073_ ( .A(_08624_ ), .B(_08625_ ), .S(fanout_net_4 ), .Z(_08626_ ) );
AND2_X1 _12074_ ( .A1(_08626_ ), .A2(_08588_ ), .ZN(_08627_ ) );
MUX2_X1 _12075_ ( .A(\u_gpr.regfile[0][0] ), .B(\u_gpr.regfile[1][0] ), .S(fanout_net_5 ), .Z(_08628_ ) );
MUX2_X1 _12076_ ( .A(\u_gpr.regfile[2][0] ), .B(\u_gpr.regfile[3][0] ), .S(fanout_net_5 ), .Z(_08629_ ) );
MUX2_X1 _12077_ ( .A(_08628_ ), .B(_08629_ ), .S(fanout_net_7 ), .Z(_08630_ ) );
AND2_X2 _12078_ ( .A1(_08630_ ), .A2(_08580_ ), .ZN(_08631_ ) );
XNOR2_X1 _12079_ ( .A(_08627_ ), .B(_08631_ ), .ZN(_08632_ ) );
MUX2_X1 _12080_ ( .A(\u_gpr.regfile[0][1] ), .B(\u_gpr.regfile[1][1] ), .S(fanout_net_5 ), .Z(_08633_ ) );
MUX2_X1 _12081_ ( .A(\u_gpr.regfile[2][1] ), .B(\u_gpr.regfile[3][1] ), .S(fanout_net_5 ), .Z(_08634_ ) );
MUX2_X1 _12082_ ( .A(_08633_ ), .B(_08634_ ), .S(fanout_net_7 ), .Z(_08635_ ) );
CLKBUF_X2 _12083_ ( .A(_08580_ ), .Z(_08636_ ) );
CLKBUF_X2 _12084_ ( .A(_08636_ ), .Z(_08637_ ) );
AND2_X1 _12085_ ( .A1(_08635_ ), .A2(_08637_ ), .ZN(_08638_ ) );
INV_X1 _12086_ ( .A(_08638_ ), .ZN(_08639_ ) );
MUX2_X1 _12087_ ( .A(\u_gpr.regfile[0][1] ), .B(\u_gpr.regfile[1][1] ), .S(fanout_net_2 ), .Z(_08640_ ) );
MUX2_X1 _12088_ ( .A(\u_gpr.regfile[2][1] ), .B(\u_gpr.regfile[3][1] ), .S(fanout_net_2 ), .Z(_08641_ ) );
MUX2_X1 _12089_ ( .A(_08640_ ), .B(_08641_ ), .S(fanout_net_4 ), .Z(_08642_ ) );
AND2_X1 _12090_ ( .A1(_08642_ ), .A2(_08611_ ), .ZN(_08643_ ) );
OR2_X1 _12091_ ( .A1(_08639_ ), .A2(_08643_ ), .ZN(_08644_ ) );
NAND2_X1 _12092_ ( .A1(_08639_ ), .A2(_08643_ ), .ZN(_08645_ ) );
NAND3_X1 _12093_ ( .A1(_08632_ ), .A2(_08644_ ), .A3(_08645_ ), .ZN(_08646_ ) );
MUX2_X1 _12094_ ( .A(\u_gpr.regfile[0][3] ), .B(\u_gpr.regfile[1][3] ), .S(fanout_net_5 ), .Z(_08647_ ) );
MUX2_X1 _12095_ ( .A(\u_gpr.regfile[2][3] ), .B(\u_gpr.regfile[3][3] ), .S(fanout_net_5 ), .Z(_08648_ ) );
MUX2_X1 _12096_ ( .A(_08647_ ), .B(_08648_ ), .S(fanout_net_7 ), .Z(_08649_ ) );
AND2_X2 _12097_ ( .A1(_08649_ ), .A2(_08580_ ), .ZN(_08650_ ) );
MUX2_X1 _12098_ ( .A(\u_gpr.regfile[0][3] ), .B(\u_gpr.regfile[1][3] ), .S(fanout_net_2 ), .Z(_08651_ ) );
MUX2_X1 _12099_ ( .A(\u_gpr.regfile[2][3] ), .B(\u_gpr.regfile[3][3] ), .S(fanout_net_2 ), .Z(_08652_ ) );
MUX2_X1 _12100_ ( .A(_08651_ ), .B(_08652_ ), .S(fanout_net_4 ), .Z(_08653_ ) );
AND2_X1 _12101_ ( .A1(_08653_ ), .A2(_08611_ ), .ZN(_08654_ ) );
XOR2_X1 _12102_ ( .A(_08650_ ), .B(_08654_ ), .Z(_08655_ ) );
MUX2_X1 _12103_ ( .A(\u_gpr.regfile[0][2] ), .B(\u_gpr.regfile[1][2] ), .S(fanout_net_5 ), .Z(_08656_ ) );
MUX2_X1 _12104_ ( .A(\u_gpr.regfile[2][2] ), .B(\u_gpr.regfile[3][2] ), .S(fanout_net_5 ), .Z(_08657_ ) );
MUX2_X1 _12105_ ( .A(_08656_ ), .B(_08657_ ), .S(fanout_net_7 ), .Z(_08658_ ) );
AND2_X2 _12106_ ( .A1(_08658_ ), .A2(_08580_ ), .ZN(_08659_ ) );
MUX2_X1 _12107_ ( .A(\u_gpr.regfile[0][2] ), .B(\u_gpr.regfile[1][2] ), .S(fanout_net_2 ), .Z(_08660_ ) );
MUX2_X1 _12108_ ( .A(\u_gpr.regfile[2][2] ), .B(\u_gpr.regfile[3][2] ), .S(fanout_net_2 ), .Z(_08661_ ) );
MUX2_X1 _12109_ ( .A(_08660_ ), .B(_08661_ ), .S(fanout_net_4 ), .Z(_08662_ ) );
NAND2_X1 _12110_ ( .A1(_08662_ ), .A2(_08588_ ), .ZN(_08663_ ) );
XNOR2_X1 _12111_ ( .A(_08659_ ), .B(_08663_ ), .ZN(_08664_ ) );
NOR4_X1 _12112_ ( .A1(_08623_ ), .A2(_08646_ ), .A3(_08655_ ), .A4(_08664_ ), .ZN(_08665_ ) );
MUX2_X1 _12113_ ( .A(\u_gpr.regfile[0][11] ), .B(\u_gpr.regfile[1][11] ), .S(fanout_net_2 ), .Z(_08666_ ) );
MUX2_X1 _12114_ ( .A(\u_gpr.regfile[2][11] ), .B(\u_gpr.regfile[3][11] ), .S(fanout_net_2 ), .Z(_08667_ ) );
MUX2_X1 _12115_ ( .A(_08666_ ), .B(_08667_ ), .S(fanout_net_4 ), .Z(_08668_ ) );
AND2_X1 _12116_ ( .A1(_08668_ ), .A2(_08589_ ), .ZN(_08669_ ) );
MUX2_X1 _12117_ ( .A(\u_gpr.regfile[0][11] ), .B(\u_gpr.regfile[1][11] ), .S(fanout_net_5 ), .Z(_08670_ ) );
MUX2_X1 _12118_ ( .A(\u_gpr.regfile[2][11] ), .B(\u_gpr.regfile[3][11] ), .S(fanout_net_5 ), .Z(_08671_ ) );
MUX2_X1 _12119_ ( .A(_08670_ ), .B(_08671_ ), .S(fanout_net_7 ), .Z(_08672_ ) );
NAND2_X1 _12120_ ( .A1(_08672_ ), .A2(_08636_ ), .ZN(_08673_ ) );
XOR2_X1 _12121_ ( .A(_08669_ ), .B(_08673_ ), .Z(_08674_ ) );
MUX2_X1 _12122_ ( .A(\u_gpr.regfile[0][8] ), .B(\u_gpr.regfile[1][8] ), .S(fanout_net_5 ), .Z(_08675_ ) );
MUX2_X1 _12123_ ( .A(\u_gpr.regfile[2][8] ), .B(\u_gpr.regfile[3][8] ), .S(fanout_net_5 ), .Z(_08676_ ) );
MUX2_X1 _12124_ ( .A(_08675_ ), .B(_08676_ ), .S(fanout_net_7 ), .Z(_08677_ ) );
AND2_X1 _12125_ ( .A1(_08677_ ), .A2(_08637_ ), .ZN(_08678_ ) );
MUX2_X1 _12126_ ( .A(\u_gpr.regfile[0][8] ), .B(\u_gpr.regfile[1][8] ), .S(fanout_net_2 ), .Z(_08679_ ) );
MUX2_X1 _12127_ ( .A(\u_gpr.regfile[2][8] ), .B(\u_gpr.regfile[3][8] ), .S(fanout_net_2 ), .Z(_08680_ ) );
MUX2_X1 _12128_ ( .A(_08679_ ), .B(_08680_ ), .S(fanout_net_4 ), .Z(_08681_ ) );
NAND2_X1 _12129_ ( .A1(_08681_ ), .A2(_08609_ ), .ZN(_08682_ ) );
XOR2_X1 _12130_ ( .A(_08678_ ), .B(_08682_ ), .Z(_08683_ ) );
MUX2_X1 _12131_ ( .A(\u_gpr.regfile[0][9] ), .B(\u_gpr.regfile[1][9] ), .S(fanout_net_5 ), .Z(_08684_ ) );
MUX2_X1 _12132_ ( .A(\u_gpr.regfile[2][9] ), .B(\u_gpr.regfile[3][9] ), .S(fanout_net_5 ), .Z(_08685_ ) );
MUX2_X1 _12133_ ( .A(_08684_ ), .B(_08685_ ), .S(fanout_net_7 ), .Z(_08686_ ) );
BUF_X2 _12134_ ( .A(_08637_ ), .Z(_08687_ ) );
NAND2_X1 _12135_ ( .A1(_08686_ ), .A2(_08687_ ), .ZN(_08688_ ) );
MUX2_X1 _12136_ ( .A(\u_gpr.regfile[0][9] ), .B(\u_gpr.regfile[1][9] ), .S(fanout_net_2 ), .Z(_08689_ ) );
MUX2_X1 _12137_ ( .A(\u_gpr.regfile[2][9] ), .B(\u_gpr.regfile[3][9] ), .S(fanout_net_2 ), .Z(_08690_ ) );
MUX2_X1 _12138_ ( .A(_08689_ ), .B(_08690_ ), .S(fanout_net_4 ), .Z(_08691_ ) );
NAND2_X1 _12139_ ( .A1(_08691_ ), .A2(_08609_ ), .ZN(_08692_ ) );
XNOR2_X1 _12140_ ( .A(_08688_ ), .B(_08692_ ), .ZN(_08693_ ) );
MUX2_X1 _12141_ ( .A(\u_gpr.regfile[0][10] ), .B(\u_gpr.regfile[1][10] ), .S(fanout_net_2 ), .Z(_08694_ ) );
MUX2_X1 _12142_ ( .A(\u_gpr.regfile[2][10] ), .B(\u_gpr.regfile[3][10] ), .S(fanout_net_2 ), .Z(_08695_ ) );
MUX2_X1 _12143_ ( .A(_08694_ ), .B(_08695_ ), .S(fanout_net_4 ), .Z(_08696_ ) );
AND2_X1 _12144_ ( .A1(_08696_ ), .A2(_08589_ ), .ZN(_08697_ ) );
INV_X1 _12145_ ( .A(fanout_net_5 ), .ZN(_08698_ ) );
OR2_X1 _12146_ ( .A1(_08698_ ), .A2(\u_gpr.regfile[3][10] ), .ZN(_08699_ ) );
OAI211_X1 _12147_ ( .A(_08699_ ), .B(fanout_net_7 ), .C1(fanout_net_5 ), .C2(\u_gpr.regfile[2][10] ), .ZN(_08700_ ) );
OR2_X1 _12148_ ( .A1(fanout_net_5 ), .A2(\u_gpr.regfile[0][10] ), .ZN(_08701_ ) );
INV_X1 _12149_ ( .A(fanout_net_7 ), .ZN(_08702_ ) );
OAI211_X1 _12150_ ( .A(_08701_ ), .B(_08702_ ), .C1(_08698_ ), .C2(\u_gpr.regfile[1][10] ), .ZN(_08703_ ) );
AOI21_X1 _12151_ ( .A(_08579_ ), .B1(_08700_ ), .B2(_08703_ ), .ZN(_08704_ ) );
XNOR2_X1 _12152_ ( .A(_08697_ ), .B(_08704_ ), .ZN(_08705_ ) );
AND4_X1 _12153_ ( .A1(_08674_ ), .A2(_08683_ ), .A3(_08693_ ), .A4(_08705_ ), .ZN(_08706_ ) );
MUX2_X1 _12154_ ( .A(\u_gpr.regfile[0][13] ), .B(\u_gpr.regfile[1][13] ), .S(fanout_net_5 ), .Z(_08707_ ) );
MUX2_X1 _12155_ ( .A(\u_gpr.regfile[2][13] ), .B(\u_gpr.regfile[3][13] ), .S(fanout_net_5 ), .Z(_08708_ ) );
MUX2_X1 _12156_ ( .A(_08707_ ), .B(_08708_ ), .S(fanout_net_7 ), .Z(_08709_ ) );
AND2_X1 _12157_ ( .A1(_08709_ ), .A2(_08636_ ), .ZN(_08710_ ) );
MUX2_X1 _12158_ ( .A(\u_gpr.regfile[0][13] ), .B(\u_gpr.regfile[1][13] ), .S(fanout_net_2 ), .Z(_08711_ ) );
MUX2_X1 _12159_ ( .A(\u_gpr.regfile[2][13] ), .B(\u_gpr.regfile[3][13] ), .S(fanout_net_2 ), .Z(_08712_ ) );
MUX2_X1 _12160_ ( .A(_08711_ ), .B(_08712_ ), .S(fanout_net_4 ), .Z(_08713_ ) );
AND2_X1 _12161_ ( .A1(_08713_ ), .A2(_08609_ ), .ZN(_08714_ ) );
XNOR2_X1 _12162_ ( .A(_08710_ ), .B(_08714_ ), .ZN(_08715_ ) );
MUX2_X1 _12163_ ( .A(\u_gpr.regfile[0][15] ), .B(\u_gpr.regfile[1][15] ), .S(fanout_net_5 ), .Z(_08716_ ) );
MUX2_X1 _12164_ ( .A(\u_gpr.regfile[2][15] ), .B(\u_gpr.regfile[3][15] ), .S(fanout_net_5 ), .Z(_08717_ ) );
MUX2_X1 _12165_ ( .A(_08716_ ), .B(_08717_ ), .S(fanout_net_7 ), .Z(_08718_ ) );
AND2_X1 _12166_ ( .A1(_08718_ ), .A2(_08687_ ), .ZN(_08719_ ) );
MUX2_X1 _12167_ ( .A(\u_gpr.regfile[0][15] ), .B(\u_gpr.regfile[1][15] ), .S(fanout_net_2 ), .Z(_08720_ ) );
MUX2_X1 _12168_ ( .A(\u_gpr.regfile[2][15] ), .B(\u_gpr.regfile[3][15] ), .S(fanout_net_2 ), .Z(_08721_ ) );
MUX2_X1 _12169_ ( .A(_08720_ ), .B(_08721_ ), .S(fanout_net_4 ), .Z(_08722_ ) );
AND2_X1 _12170_ ( .A1(_08722_ ), .A2(_08609_ ), .ZN(_08723_ ) );
XNOR2_X1 _12171_ ( .A(_08719_ ), .B(_08723_ ), .ZN(_08724_ ) );
MUX2_X1 _12172_ ( .A(\u_gpr.regfile[0][12] ), .B(\u_gpr.regfile[1][12] ), .S(fanout_net_2 ), .Z(_08725_ ) );
MUX2_X1 _12173_ ( .A(\u_gpr.regfile[2][12] ), .B(\u_gpr.regfile[3][12] ), .S(fanout_net_3 ), .Z(_08726_ ) );
MUX2_X1 _12174_ ( .A(_08725_ ), .B(_08726_ ), .S(fanout_net_4 ), .Z(_08727_ ) );
AND2_X1 _12175_ ( .A1(_08727_ ), .A2(_08609_ ), .ZN(_08728_ ) );
MUX2_X1 _12176_ ( .A(\u_gpr.regfile[0][12] ), .B(\u_gpr.regfile[1][12] ), .S(fanout_net_6 ), .Z(_08729_ ) );
MUX2_X1 _12177_ ( .A(\u_gpr.regfile[2][12] ), .B(\u_gpr.regfile[3][12] ), .S(fanout_net_6 ), .Z(_08730_ ) );
MUX2_X1 _12178_ ( .A(_08729_ ), .B(_08730_ ), .S(fanout_net_7 ), .Z(_08731_ ) );
AND2_X1 _12179_ ( .A1(_08731_ ), .A2(_08636_ ), .ZN(_08732_ ) );
XNOR2_X1 _12180_ ( .A(_08728_ ), .B(_08732_ ), .ZN(_08733_ ) );
MUX2_X1 _12181_ ( .A(\u_gpr.regfile[0][14] ), .B(\u_gpr.regfile[1][14] ), .S(fanout_net_3 ), .Z(_08734_ ) );
MUX2_X1 _12182_ ( .A(\u_gpr.regfile[2][14] ), .B(\u_gpr.regfile[3][14] ), .S(fanout_net_3 ), .Z(_08735_ ) );
MUX2_X1 _12183_ ( .A(_08734_ ), .B(_08735_ ), .S(fanout_net_4 ), .Z(_08736_ ) );
AND2_X1 _12184_ ( .A1(_08736_ ), .A2(_08589_ ), .ZN(_08737_ ) );
MUX2_X1 _12185_ ( .A(\u_gpr.regfile[0][14] ), .B(\u_gpr.regfile[1][14] ), .S(fanout_net_6 ), .Z(_08738_ ) );
MUX2_X1 _12186_ ( .A(\u_gpr.regfile[2][14] ), .B(\u_gpr.regfile[3][14] ), .S(fanout_net_6 ), .Z(_08739_ ) );
MUX2_X1 _12187_ ( .A(_08738_ ), .B(_08739_ ), .S(fanout_net_7 ), .Z(_08740_ ) );
AND2_X1 _12188_ ( .A1(_08740_ ), .A2(_08636_ ), .ZN(_08741_ ) );
XNOR2_X1 _12189_ ( .A(_08737_ ), .B(_08741_ ), .ZN(_08742_ ) );
AND4_X1 _12190_ ( .A1(_08715_ ), .A2(_08724_ ), .A3(_08733_ ), .A4(_08742_ ), .ZN(_08743_ ) );
NAND3_X1 _12191_ ( .A1(_08665_ ), .A2(_08706_ ), .A3(_08743_ ), .ZN(_08744_ ) );
MUX2_X1 _12192_ ( .A(\u_gpr.regfile[0][19] ), .B(\u_gpr.regfile[1][19] ), .S(fanout_net_6 ), .Z(_08745_ ) );
MUX2_X1 _12193_ ( .A(\u_gpr.regfile[2][19] ), .B(\u_gpr.regfile[3][19] ), .S(fanout_net_6 ), .Z(_08746_ ) );
MUX2_X1 _12194_ ( .A(_08745_ ), .B(_08746_ ), .S(fanout_net_7 ), .Z(_08747_ ) );
AND2_X1 _12195_ ( .A1(_08747_ ), .A2(_08636_ ), .ZN(_08748_ ) );
MUX2_X1 _12196_ ( .A(\u_gpr.regfile[0][19] ), .B(\u_gpr.regfile[1][19] ), .S(fanout_net_3 ), .Z(_08749_ ) );
MUX2_X1 _12197_ ( .A(\u_gpr.regfile[2][19] ), .B(\u_gpr.regfile[3][19] ), .S(fanout_net_3 ), .Z(_08750_ ) );
MUX2_X1 _12198_ ( .A(_08749_ ), .B(_08750_ ), .S(fanout_net_4 ), .Z(_08751_ ) );
AND2_X1 _12199_ ( .A1(_08751_ ), .A2(_08609_ ), .ZN(_08752_ ) );
XNOR2_X1 _12200_ ( .A(_08748_ ), .B(_08752_ ), .ZN(_08753_ ) );
MUX2_X1 _12201_ ( .A(\u_gpr.regfile[0][18] ), .B(\u_gpr.regfile[1][18] ), .S(fanout_net_6 ), .Z(_08754_ ) );
MUX2_X1 _12202_ ( .A(\u_gpr.regfile[2][18] ), .B(\u_gpr.regfile[3][18] ), .S(fanout_net_6 ), .Z(_08755_ ) );
MUX2_X1 _12203_ ( .A(_08754_ ), .B(_08755_ ), .S(fanout_net_7 ), .Z(_08756_ ) );
NAND2_X1 _12204_ ( .A1(_08756_ ), .A2(_08687_ ), .ZN(_08757_ ) );
MUX2_X1 _12205_ ( .A(\u_gpr.regfile[0][18] ), .B(\u_gpr.regfile[1][18] ), .S(fanout_net_3 ), .Z(_08758_ ) );
MUX2_X1 _12206_ ( .A(\u_gpr.regfile[2][18] ), .B(\u_gpr.regfile[3][18] ), .S(fanout_net_3 ), .Z(_08759_ ) );
MUX2_X1 _12207_ ( .A(_08758_ ), .B(_08759_ ), .S(fanout_net_4 ), .Z(_08760_ ) );
NAND3_X1 _12208_ ( .A1(_08757_ ), .A2(_08611_ ), .A3(_08760_ ), .ZN(_08761_ ) );
AND2_X1 _12209_ ( .A1(_08760_ ), .A2(_08609_ ), .ZN(_08762_ ) );
OR2_X1 _12210_ ( .A1(_08762_ ), .A2(_08757_ ), .ZN(_08763_ ) );
AND3_X1 _12211_ ( .A1(_08753_ ), .A2(_08761_ ), .A3(_08763_ ), .ZN(_08764_ ) );
MUX2_X1 _12212_ ( .A(\u_gpr.regfile[0][16] ), .B(\u_gpr.regfile[1][16] ), .S(fanout_net_6 ), .Z(_08765_ ) );
MUX2_X1 _12213_ ( .A(\u_gpr.regfile[2][16] ), .B(\u_gpr.regfile[3][16] ), .S(fanout_net_6 ), .Z(_08766_ ) );
MUX2_X1 _12214_ ( .A(_08765_ ), .B(_08766_ ), .S(fanout_net_7 ), .Z(_08767_ ) );
AND2_X1 _12215_ ( .A1(_08767_ ), .A2(_08636_ ), .ZN(_08768_ ) );
MUX2_X1 _12216_ ( .A(\u_gpr.regfile[0][16] ), .B(\u_gpr.regfile[1][16] ), .S(fanout_net_3 ), .Z(_08769_ ) );
MUX2_X1 _12217_ ( .A(\u_gpr.regfile[2][16] ), .B(\u_gpr.regfile[3][16] ), .S(fanout_net_3 ), .Z(_08770_ ) );
MUX2_X1 _12218_ ( .A(_08769_ ), .B(_08770_ ), .S(fanout_net_4 ), .Z(_08771_ ) );
AND2_X1 _12219_ ( .A1(_08771_ ), .A2(_08609_ ), .ZN(_08772_ ) );
XNOR2_X1 _12220_ ( .A(_08768_ ), .B(_08772_ ), .ZN(_08773_ ) );
MUX2_X1 _12221_ ( .A(\u_gpr.regfile[0][17] ), .B(\u_gpr.regfile[1][17] ), .S(fanout_net_6 ), .Z(_08774_ ) );
MUX2_X1 _12222_ ( .A(\u_gpr.regfile[2][17] ), .B(\u_gpr.regfile[3][17] ), .S(fanout_net_6 ), .Z(_08775_ ) );
MUX2_X1 _12223_ ( .A(_08774_ ), .B(_08775_ ), .S(fanout_net_7 ), .Z(_08776_ ) );
MUX2_X1 _12224_ ( .A(\u_gpr.regfile[0][17] ), .B(\u_gpr.regfile[1][17] ), .S(fanout_net_3 ), .Z(_08777_ ) );
MUX2_X1 _12225_ ( .A(\u_gpr.regfile[2][17] ), .B(\u_gpr.regfile[3][17] ), .S(fanout_net_3 ), .Z(_08778_ ) );
MUX2_X1 _12226_ ( .A(_08777_ ), .B(_08778_ ), .S(fanout_net_4 ), .Z(_08779_ ) );
AND4_X1 _12227_ ( .A1(_08687_ ), .A2(_08776_ ), .A3(_08779_ ), .A4(_08611_ ), .ZN(_08780_ ) );
AOI22_X1 _12228_ ( .A1(_08687_ ), .A2(_08776_ ), .B1(_08779_ ), .B2(_08611_ ), .ZN(_08781_ ) );
OAI211_X1 _12229_ ( .A(_08764_ ), .B(_08773_ ), .C1(_08780_ ), .C2(_08781_ ), .ZN(_08782_ ) );
MUX2_X1 _12230_ ( .A(\u_gpr.regfile[0][20] ), .B(\u_gpr.regfile[1][20] ), .S(fanout_net_3 ), .Z(_08783_ ) );
MUX2_X1 _12231_ ( .A(\u_gpr.regfile[2][20] ), .B(\u_gpr.regfile[3][20] ), .S(fanout_net_3 ), .Z(_08784_ ) );
MUX2_X1 _12232_ ( .A(_08783_ ), .B(_08784_ ), .S(fanout_net_4 ), .Z(_08785_ ) );
AND2_X1 _12233_ ( .A1(_08785_ ), .A2(_08610_ ), .ZN(_08786_ ) );
MUX2_X1 _12234_ ( .A(\u_gpr.regfile[0][20] ), .B(\u_gpr.regfile[1][20] ), .S(fanout_net_6 ), .Z(_08787_ ) );
MUX2_X1 _12235_ ( .A(\u_gpr.regfile[2][20] ), .B(\u_gpr.regfile[3][20] ), .S(fanout_net_6 ), .Z(_08788_ ) );
MUX2_X1 _12236_ ( .A(_08787_ ), .B(_08788_ ), .S(fanout_net_7 ), .Z(_08789_ ) );
NAND2_X1 _12237_ ( .A1(_08789_ ), .A2(_08687_ ), .ZN(_08790_ ) );
XOR2_X1 _12238_ ( .A(_08786_ ), .B(_08790_ ), .Z(_08791_ ) );
MUX2_X1 _12239_ ( .A(\u_gpr.regfile[0][21] ), .B(\u_gpr.regfile[1][21] ), .S(fanout_net_6 ), .Z(_08792_ ) );
MUX2_X1 _12240_ ( .A(\u_gpr.regfile[2][21] ), .B(\u_gpr.regfile[3][21] ), .S(fanout_net_6 ), .Z(_08793_ ) );
MUX2_X1 _12241_ ( .A(_08792_ ), .B(_08793_ ), .S(fanout_net_7 ), .Z(_08794_ ) );
AND2_X1 _12242_ ( .A1(_08794_ ), .A2(_08637_ ), .ZN(_08795_ ) );
MUX2_X1 _12243_ ( .A(\u_gpr.regfile[0][21] ), .B(\u_gpr.regfile[1][21] ), .S(fanout_net_3 ), .Z(_08796_ ) );
MUX2_X1 _12244_ ( .A(\u_gpr.regfile[2][21] ), .B(\u_gpr.regfile[3][21] ), .S(fanout_net_3 ), .Z(_08797_ ) );
MUX2_X1 _12245_ ( .A(_08796_ ), .B(_08797_ ), .S(fanout_net_4 ), .Z(_08798_ ) );
AND2_X1 _12246_ ( .A1(_08798_ ), .A2(_08609_ ), .ZN(_08799_ ) );
XNOR2_X1 _12247_ ( .A(_08795_ ), .B(_08799_ ), .ZN(_08800_ ) );
MUX2_X1 _12248_ ( .A(\u_gpr.regfile[0][23] ), .B(\u_gpr.regfile[1][23] ), .S(fanout_net_6 ), .Z(_08801_ ) );
MUX2_X1 _12249_ ( .A(\u_gpr.regfile[2][23] ), .B(\u_gpr.regfile[3][23] ), .S(fanout_net_6 ), .Z(_08802_ ) );
MUX2_X1 _12250_ ( .A(_08801_ ), .B(_08802_ ), .S(fanout_net_7 ), .Z(_08803_ ) );
AND2_X1 _12251_ ( .A1(_08803_ ), .A2(_08637_ ), .ZN(_08804_ ) );
MUX2_X1 _12252_ ( .A(\u_gpr.regfile[0][23] ), .B(\u_gpr.regfile[1][23] ), .S(fanout_net_3 ), .Z(_08805_ ) );
MUX2_X1 _12253_ ( .A(\u_gpr.regfile[2][23] ), .B(\u_gpr.regfile[3][23] ), .S(fanout_net_3 ), .Z(_08806_ ) );
MUX2_X1 _12254_ ( .A(_08805_ ), .B(_08806_ ), .S(fanout_net_4 ), .Z(_08807_ ) );
AND2_X1 _12255_ ( .A1(_08807_ ), .A2(_08610_ ), .ZN(_08808_ ) );
XNOR2_X1 _12256_ ( .A(_08804_ ), .B(_08808_ ), .ZN(_08809_ ) );
MUX2_X1 _12257_ ( .A(\u_gpr.regfile[0][22] ), .B(\u_gpr.regfile[1][22] ), .S(fanout_net_3 ), .Z(_08810_ ) );
MUX2_X1 _12258_ ( .A(\u_gpr.regfile[2][22] ), .B(\u_gpr.regfile[3][22] ), .S(fanout_net_3 ), .Z(_08811_ ) );
MUX2_X1 _12259_ ( .A(_08810_ ), .B(_08811_ ), .S(fanout_net_4 ), .Z(_08812_ ) );
AND2_X1 _12260_ ( .A1(_08812_ ), .A2(_08610_ ), .ZN(_08813_ ) );
OR2_X1 _12261_ ( .A1(_08698_ ), .A2(\u_gpr.regfile[3][22] ), .ZN(_08814_ ) );
OAI211_X1 _12262_ ( .A(_08814_ ), .B(fanout_net_7 ), .C1(fanout_net_6 ), .C2(\u_gpr.regfile[2][22] ), .ZN(_08815_ ) );
OR2_X1 _12263_ ( .A1(fanout_net_6 ), .A2(\u_gpr.regfile[0][22] ), .ZN(_08816_ ) );
OAI211_X1 _12264_ ( .A(_08816_ ), .B(_08702_ ), .C1(_08698_ ), .C2(\u_gpr.regfile[1][22] ), .ZN(_08817_ ) );
AOI21_X1 _12265_ ( .A(_08579_ ), .B1(_08815_ ), .B2(_08817_ ), .ZN(_08818_ ) );
XNOR2_X1 _12266_ ( .A(_08813_ ), .B(_08818_ ), .ZN(_08819_ ) );
NAND4_X1 _12267_ ( .A1(_08791_ ), .A2(_08800_ ), .A3(_08809_ ), .A4(_08819_ ), .ZN(_08820_ ) );
MUX2_X1 _12268_ ( .A(\u_gpr.regfile[0][29] ), .B(\u_gpr.regfile[1][29] ), .S(fanout_net_6 ), .Z(_08821_ ) );
MUX2_X1 _12269_ ( .A(\u_gpr.regfile[2][29] ), .B(\u_gpr.regfile[3][29] ), .S(fanout_net_6 ), .Z(_08822_ ) );
MUX2_X1 _12270_ ( .A(_08821_ ), .B(_08822_ ), .S(fanout_net_7 ), .Z(_08823_ ) );
AND2_X1 _12271_ ( .A1(_08823_ ), .A2(_08637_ ), .ZN(_08824_ ) );
MUX2_X1 _12272_ ( .A(\u_gpr.regfile[0][29] ), .B(\u_gpr.regfile[1][29] ), .S(fanout_net_3 ), .Z(_08825_ ) );
MUX2_X1 _12273_ ( .A(\u_gpr.regfile[2][29] ), .B(\u_gpr.regfile[3][29] ), .S(fanout_net_3 ), .Z(_08826_ ) );
MUX2_X1 _12274_ ( .A(_08825_ ), .B(_08826_ ), .S(fanout_net_4 ), .Z(_08827_ ) );
NAND2_X1 _12275_ ( .A1(_08827_ ), .A2(_08611_ ), .ZN(_08828_ ) );
XOR2_X1 _12276_ ( .A(_08824_ ), .B(_08828_ ), .Z(_08829_ ) );
MUX2_X1 _12277_ ( .A(\u_gpr.regfile[0][31] ), .B(\u_gpr.regfile[1][31] ), .S(fanout_net_3 ), .Z(_08830_ ) );
MUX2_X1 _12278_ ( .A(\u_gpr.regfile[2][31] ), .B(\u_gpr.regfile[3][31] ), .S(fanout_net_3 ), .Z(_08831_ ) );
MUX2_X1 _12279_ ( .A(_08830_ ), .B(_08831_ ), .S(fanout_net_4 ), .Z(_08832_ ) );
AND2_X1 _12280_ ( .A1(_08832_ ), .A2(_08610_ ), .ZN(_08833_ ) );
MUX2_X1 _12281_ ( .A(\u_gpr.regfile[0][31] ), .B(\u_gpr.regfile[1][31] ), .S(fanout_net_6 ), .Z(_08834_ ) );
MUX2_X1 _12282_ ( .A(\u_gpr.regfile[2][31] ), .B(\u_gpr.regfile[3][31] ), .S(fanout_net_6 ), .Z(_08835_ ) );
MUX2_X1 _12283_ ( .A(_08834_ ), .B(_08835_ ), .S(fanout_net_7 ), .Z(_08836_ ) );
NAND2_X1 _12284_ ( .A1(_08836_ ), .A2(_08687_ ), .ZN(_08837_ ) );
XOR2_X1 _12285_ ( .A(_08833_ ), .B(_08837_ ), .Z(_08838_ ) );
MUX2_X1 _12286_ ( .A(\u_gpr.regfile[0][28] ), .B(\u_gpr.regfile[1][28] ), .S(fanout_net_3 ), .Z(_08839_ ) );
MUX2_X1 _12287_ ( .A(\u_gpr.regfile[2][28] ), .B(\u_gpr.regfile[3][28] ), .S(fanout_net_3 ), .Z(_08840_ ) );
MUX2_X1 _12288_ ( .A(_08839_ ), .B(_08840_ ), .S(fanout_net_4 ), .Z(_08841_ ) );
AND2_X1 _12289_ ( .A1(_08841_ ), .A2(_08610_ ), .ZN(_08842_ ) );
MUX2_X1 _12290_ ( .A(\u_gpr.regfile[0][28] ), .B(\u_gpr.regfile[1][28] ), .S(fanout_net_6 ), .Z(_08843_ ) );
MUX2_X1 _12291_ ( .A(\u_gpr.regfile[2][28] ), .B(\u_gpr.regfile[3][28] ), .S(fanout_net_6 ), .Z(_08844_ ) );
MUX2_X1 _12292_ ( .A(_08843_ ), .B(_08844_ ), .S(fanout_net_7 ), .Z(_08845_ ) );
AND2_X1 _12293_ ( .A1(_08845_ ), .A2(_08637_ ), .ZN(_08846_ ) );
XNOR2_X1 _12294_ ( .A(_08842_ ), .B(_08846_ ), .ZN(_08847_ ) );
MUX2_X1 _12295_ ( .A(\u_gpr.regfile[0][30] ), .B(\u_gpr.regfile[1][30] ), .S(fanout_net_3 ), .Z(_08848_ ) );
MUX2_X1 _12296_ ( .A(\u_gpr.regfile[2][30] ), .B(\u_gpr.regfile[3][30] ), .S(fanout_net_3 ), .Z(_08849_ ) );
MUX2_X1 _12297_ ( .A(_08848_ ), .B(_08849_ ), .S(fanout_net_4 ), .Z(_08850_ ) );
NAND2_X1 _12298_ ( .A1(_08850_ ), .A2(_08611_ ), .ZN(_08851_ ) );
OR2_X1 _12299_ ( .A1(_08698_ ), .A2(\u_gpr.regfile[1][30] ), .ZN(_08852_ ) );
OAI211_X1 _12300_ ( .A(_08852_ ), .B(_08702_ ), .C1(fanout_net_6 ), .C2(\u_gpr.regfile[0][30] ), .ZN(_08853_ ) );
OR2_X1 _12301_ ( .A1(fanout_net_6 ), .A2(\u_gpr.regfile[2][30] ), .ZN(_08854_ ) );
OAI211_X1 _12302_ ( .A(_08854_ ), .B(fanout_net_7 ), .C1(_08698_ ), .C2(\u_gpr.regfile[3][30] ), .ZN(_08855_ ) );
AOI21_X1 _12303_ ( .A(_08579_ ), .B1(_08853_ ), .B2(_08855_ ), .ZN(_08856_ ) );
XOR2_X1 _12304_ ( .A(_08851_ ), .B(_08856_ ), .Z(_08857_ ) );
AND4_X1 _12305_ ( .A1(_08829_ ), .A2(_08838_ ), .A3(_08847_ ), .A4(_08857_ ), .ZN(_08858_ ) );
MUX2_X1 _12306_ ( .A(\u_gpr.regfile[0][25] ), .B(\u_gpr.regfile[1][25] ), .S(fanout_net_6 ), .Z(_08859_ ) );
MUX2_X1 _12307_ ( .A(\u_gpr.regfile[2][25] ), .B(\u_gpr.regfile[3][25] ), .S(fanout_net_6 ), .Z(_08860_ ) );
MUX2_X1 _12308_ ( .A(_08859_ ), .B(_08860_ ), .S(\ifu_rdata[21] ), .Z(_08861_ ) );
AND2_X1 _12309_ ( .A1(_08861_ ), .A2(_08637_ ), .ZN(_08862_ ) );
MUX2_X1 _12310_ ( .A(\u_gpr.regfile[0][25] ), .B(\u_gpr.regfile[1][25] ), .S(fanout_net_3 ), .Z(_08863_ ) );
MUX2_X1 _12311_ ( .A(\u_gpr.regfile[2][25] ), .B(\u_gpr.regfile[3][25] ), .S(fanout_net_3 ), .Z(_08864_ ) );
MUX2_X1 _12312_ ( .A(_08863_ ), .B(_08864_ ), .S(fanout_net_4 ), .Z(_08865_ ) );
AND2_X1 _12313_ ( .A1(_08865_ ), .A2(_08610_ ), .ZN(_08866_ ) );
XNOR2_X1 _12314_ ( .A(_08862_ ), .B(_08866_ ), .ZN(_08867_ ) );
MUX2_X1 _12315_ ( .A(\u_gpr.regfile[0][24] ), .B(\u_gpr.regfile[1][24] ), .S(fanout_net_3 ), .Z(_08868_ ) );
MUX2_X1 _12316_ ( .A(\u_gpr.regfile[2][24] ), .B(\u_gpr.regfile[3][24] ), .S(\ifu_rdata[15] ), .Z(_08869_ ) );
MUX2_X1 _12317_ ( .A(_08868_ ), .B(_08869_ ), .S(\ifu_rdata[16] ), .Z(_08870_ ) );
AND2_X1 _12318_ ( .A1(_08870_ ), .A2(_08610_ ), .ZN(_08871_ ) );
OR2_X1 _12319_ ( .A1(_08698_ ), .A2(\u_gpr.regfile[3][24] ), .ZN(_08872_ ) );
OAI211_X1 _12320_ ( .A(_08872_ ), .B(\ifu_rdata[21] ), .C1(\ifu_rdata[20] ), .C2(\u_gpr.regfile[2][24] ), .ZN(_08873_ ) );
OR2_X1 _12321_ ( .A1(_08698_ ), .A2(\u_gpr.regfile[1][24] ), .ZN(_08874_ ) );
OAI211_X1 _12322_ ( .A(_08874_ ), .B(_08702_ ), .C1(\ifu_rdata[20] ), .C2(\u_gpr.regfile[0][24] ), .ZN(_08875_ ) );
AOI21_X1 _12323_ ( .A(_08579_ ), .B1(_08873_ ), .B2(_08875_ ), .ZN(_08876_ ) );
XNOR2_X1 _12324_ ( .A(_08871_ ), .B(_08876_ ), .ZN(_08877_ ) );
MUX2_X1 _12325_ ( .A(\u_gpr.regfile[0][27] ), .B(\u_gpr.regfile[1][27] ), .S(\ifu_rdata[15] ), .Z(_08878_ ) );
MUX2_X1 _12326_ ( .A(\u_gpr.regfile[2][27] ), .B(\u_gpr.regfile[3][27] ), .S(\ifu_rdata[15] ), .Z(_08879_ ) );
MUX2_X1 _12327_ ( .A(_08878_ ), .B(_08879_ ), .S(\ifu_rdata[16] ), .Z(_08880_ ) );
AND2_X1 _12328_ ( .A1(_08880_ ), .A2(_08610_ ), .ZN(_08881_ ) );
MUX2_X1 _12329_ ( .A(\u_gpr.regfile[0][27] ), .B(\u_gpr.regfile[1][27] ), .S(\ifu_rdata[20] ), .Z(_08882_ ) );
MUX2_X1 _12330_ ( .A(\u_gpr.regfile[2][27] ), .B(\u_gpr.regfile[3][27] ), .S(\ifu_rdata[20] ), .Z(_08883_ ) );
MUX2_X1 _12331_ ( .A(_08882_ ), .B(_08883_ ), .S(\ifu_rdata[21] ), .Z(_08884_ ) );
NAND2_X1 _12332_ ( .A1(_08884_ ), .A2(_08687_ ), .ZN(_08885_ ) );
XNOR2_X1 _12333_ ( .A(_08881_ ), .B(_08885_ ), .ZN(_08886_ ) );
MUX2_X1 _12334_ ( .A(\u_gpr.regfile[0][26] ), .B(\u_gpr.regfile[1][26] ), .S(\ifu_rdata[20] ), .Z(_08887_ ) );
MUX2_X1 _12335_ ( .A(\u_gpr.regfile[2][26] ), .B(\u_gpr.regfile[3][26] ), .S(\ifu_rdata[20] ), .Z(_08888_ ) );
MUX2_X1 _12336_ ( .A(_08887_ ), .B(_08888_ ), .S(\ifu_rdata[21] ), .Z(_08889_ ) );
AND2_X1 _12337_ ( .A1(_08889_ ), .A2(_08687_ ), .ZN(_08890_ ) );
INV_X1 _12338_ ( .A(_08890_ ), .ZN(_08891_ ) );
MUX2_X1 _12339_ ( .A(\u_gpr.regfile[0][26] ), .B(\u_gpr.regfile[1][26] ), .S(\ifu_rdata[15] ), .Z(_08892_ ) );
MUX2_X1 _12340_ ( .A(\u_gpr.regfile[2][26] ), .B(\u_gpr.regfile[3][26] ), .S(\ifu_rdata[15] ), .Z(_08893_ ) );
MUX2_X1 _12341_ ( .A(_08892_ ), .B(_08893_ ), .S(\ifu_rdata[16] ), .Z(_08894_ ) );
AND2_X1 _12342_ ( .A1(_08894_ ), .A2(_08610_ ), .ZN(_08895_ ) );
AND2_X1 _12343_ ( .A1(_08891_ ), .A2(_08895_ ), .ZN(_08896_ ) );
NOR2_X1 _12344_ ( .A1(_08891_ ), .A2(_08895_ ), .ZN(_08897_ ) );
NOR3_X1 _12345_ ( .A1(_08886_ ), .A2(_08896_ ), .A3(_08897_ ), .ZN(_08898_ ) );
NAND4_X1 _12346_ ( .A1(_08858_ ), .A2(_08867_ ), .A3(_08877_ ), .A4(_08898_ ), .ZN(_08899_ ) );
NOR4_X1 _12347_ ( .A1(_08744_ ), .A2(_08782_ ), .A3(_08820_ ), .A4(_08899_ ), .ZN(_08900_ ) );
INV_X16 _12348_ ( .A(\ifu_rdata[0] ), .ZN(_08901_ ) );
NOR2_X2 _12349_ ( .A1(_08901_ ), .A2(\ifu_rdata[2] ), .ZN(_08902_ ) );
INV_X32 _12350_ ( .A(\ifu_rdata[5] ), .ZN(_08903_ ) );
NOR3_X4 _12351_ ( .A1(_08903_ ), .A2(\ifu_rdata[4] ), .A3(alu_result_out_$_XNOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B_$_OR__Y_B_$_NOR__Y_A_$_XOR__Y_B_$_OR__Y_A_$_OR__Y_B ), .ZN(_08904_ ) );
BUF_X2 _12352_ ( .A(_08904_ ), .Z(_08905_ ) );
NAND3_X1 _12353_ ( .A1(_08900_ ), .A2(_08902_ ), .A3(_08905_ ), .ZN(_08906_ ) );
AND2_X4 _12354_ ( .A1(_08904_ ), .A2(\ifu_rdata[0] ), .ZN(_08907_ ) );
AND2_X4 _12355_ ( .A1(_08907_ ), .A2(\ifu_rdata[2] ), .ZN(_08908_ ) );
INV_X4 _12356_ ( .A(_08908_ ), .ZN(_08909_ ) );
INV_X1 _12357_ ( .A(\ifu_rdata[4] ), .ZN(_08910_ ) );
OR3_X2 _12358_ ( .A1(_08910_ ), .A2(_08903_ ), .A3(alu_result_out_$_XNOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B_$_OR__Y_B_$_NOR__Y_A_$_XOR__Y_B_$_OR__Y_A_$_OR__Y_B ), .ZN(_08911_ ) );
INV_X1 _12359_ ( .A(_08902_ ), .ZN(_08912_ ) );
NOR2_X4 _12360_ ( .A1(_08911_ ), .A2(_08912_ ), .ZN(_08913_ ) );
AND2_X1 _12361_ ( .A1(_08902_ ), .A2(_08903_ ), .ZN(_08914_ ) );
NOR2_X4 _12362_ ( .A1(_08913_ ), .A2(_08914_ ), .ZN(_08915_ ) );
AOI21_X4 _12363_ ( .A(\u_ifu.jump_en_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_NOR__Y_A_$_OR__Y_B ), .B1(_08909_ ), .B2(_08915_ ), .ZN(_08916_ ) );
NOR2_X1 _12364_ ( .A1(_08903_ ), .A2(\ifu_rdata[4] ), .ZN(_08917_ ) );
AND3_X1 _12365_ ( .A1(_08902_ ), .A2(_08917_ ), .A3(\ifu_rdata[8] ), .ZN(_08918_ ) );
NOR2_X1 _12366_ ( .A1(_08916_ ), .A2(_08918_ ), .ZN(_08919_ ) );
AND2_X1 _12367_ ( .A1(_08902_ ), .A2(_08917_ ), .ZN(_08920_ ) );
BUF_X4 _12368_ ( .A(_08907_ ), .Z(_08921_ ) );
INV_X4 _12369_ ( .A(_08921_ ), .ZN(_08922_ ) );
NAND4_X1 _12370_ ( .A1(_08915_ ), .A2(\ifu_rdata[7] ), .A3(_08920_ ), .A4(_08922_ ), .ZN(_08923_ ) );
INV_X1 _12371_ ( .A(alu_result_out_$_XNOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B_$_ORNOT__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_08924_ ) );
OAI21_X1 _12372_ ( .A(_08924_ ), .B1(_08913_ ), .B2(_08914_ ), .ZN(_08925_ ) );
AND2_X1 _12373_ ( .A1(_08923_ ), .A2(_08925_ ), .ZN(_08926_ ) );
NAND3_X1 _12374_ ( .A1(_08919_ ), .A2(_08913_ ), .A3(_08926_ ), .ZN(_08927_ ) );
BUF_X2 _12375_ ( .A(_08909_ ), .Z(_08928_ ) );
AND2_X1 _12376_ ( .A1(_08927_ ), .A2(_08928_ ), .ZN(_08929_ ) );
AND2_X2 _12377_ ( .A1(_08906_ ), .A2(_08929_ ), .ZN(_08930_ ) );
INV_X1 _12378_ ( .A(_08930_ ), .ZN(_08931_ ) );
INV_X1 _12379_ ( .A(dnpc_$_NOT__Y_3_A_$_MUX__Y_A_$_XOR__Y_B ), .ZN(_08932_ ) );
MUX2_X1 _12380_ ( .A(_08932_ ), .B(_08621_ ), .S(_08922_ ), .Z(_08933_ ) );
AOI21_X4 _12381_ ( .A(_08920_ ), .B1(_08907_ ), .B2(\ifu_rdata[2] ), .ZN(_08934_ ) );
AND2_X2 _12382_ ( .A1(_08915_ ), .A2(_08934_ ), .ZN(_08935_ ) );
AND2_X1 _12383_ ( .A1(_08935_ ), .A2(_08617_ ), .ZN(_08936_ ) );
XOR2_X1 _12384_ ( .A(_08933_ ), .B(_08936_ ), .Z(_08937_ ) );
NAND2_X1 _12385_ ( .A1(_08935_ ), .A2(_08650_ ), .ZN(_08938_ ) );
NAND3_X1 _12386_ ( .A1(_08653_ ), .A2(_08589_ ), .A3(_08922_ ), .ZN(_08939_ ) );
NAND3_X1 _12387_ ( .A1(_08904_ ), .A2(\ifu_rdata[0] ), .A3(\pc_out[3] ), .ZN(_08940_ ) );
NAND2_X1 _12388_ ( .A1(_08939_ ), .A2(_08940_ ), .ZN(_08941_ ) );
XNOR2_X1 _12389_ ( .A(_08938_ ), .B(_08941_ ), .ZN(_08942_ ) );
INV_X1 _12390_ ( .A(_08942_ ), .ZN(_08943_ ) );
BUF_X4 _12391_ ( .A(_08915_ ), .Z(_08944_ ) );
NAND4_X1 _12392_ ( .A1(_08944_ ), .A2(_08635_ ), .A3(_08580_ ), .A4(_08934_ ), .ZN(_08945_ ) );
NAND2_X2 _12393_ ( .A1(_08919_ ), .A2(_08945_ ), .ZN(_08946_ ) );
AOI21_X1 _12394_ ( .A(_08921_ ), .B1(_08642_ ), .B2(_08588_ ), .ZN(_08947_ ) );
AND3_X1 _12395_ ( .A1(_08904_ ), .A2(\ifu_rdata[0] ), .A3(\u_gpr.gpr_wdata_$_ANDNOT__Y_30_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_08948_ ) );
NOR2_X4 _12396_ ( .A1(_08947_ ), .A2(_08948_ ), .ZN(_08949_ ) );
NAND2_X1 _12397_ ( .A1(_08946_ ), .A2(_08949_ ), .ZN(_08950_ ) );
XNOR2_X2 _12398_ ( .A(_08946_ ), .B(_08949_ ), .ZN(_08951_ ) );
INV_X1 _12399_ ( .A(_08631_ ), .ZN(_08952_ ) );
INV_X1 _12400_ ( .A(_08935_ ), .ZN(_08953_ ) );
OAI21_X1 _12401_ ( .A(_08926_ ), .B1(_08952_ ), .B2(_08953_ ), .ZN(_08954_ ) );
MUX2_X1 _12402_ ( .A(\pc_out[0] ), .B(_08627_ ), .S(_08922_ ), .Z(_08955_ ) );
NAND2_X1 _12403_ ( .A1(_08954_ ), .A2(_08955_ ), .ZN(_08956_ ) );
OAI21_X2 _12404_ ( .A(_08950_ ), .B1(_08951_ ), .B2(_08956_ ), .ZN(_08957_ ) );
NAND4_X1 _12405_ ( .A1(_08944_ ), .A2(\ifu_rdata[16] ), .A3(_08920_ ), .A4(_08922_ ), .ZN(_08958_ ) );
INV_X1 _12406_ ( .A(alu_result_out_$_XNOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B_$_OR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_08959_ ) );
NAND3_X1 _12407_ ( .A1(_08904_ ), .A2(_08959_ ), .A3(_08902_ ), .ZN(_08960_ ) );
AND2_X1 _12408_ ( .A1(_08958_ ), .A2(_08960_ ), .ZN(_08961_ ) );
INV_X1 _12409_ ( .A(_08659_ ), .ZN(_08962_ ) );
OAI21_X1 _12410_ ( .A(_08961_ ), .B1(_08962_ ), .B2(_08953_ ), .ZN(_08963_ ) );
INV_X1 _12411_ ( .A(dnpc_$_MUX__Y_22_A ), .ZN(_08964_ ) );
NAND3_X1 _12412_ ( .A1(_08904_ ), .A2(\ifu_rdata[0] ), .A3(_08964_ ), .ZN(_08965_ ) );
OAI21_X1 _12413_ ( .A(_08965_ ), .B1(_08663_ ), .B2(_08921_ ), .ZN(_08966_ ) );
XOR2_X1 _12414_ ( .A(_08963_ ), .B(_08966_ ), .Z(_08967_ ) );
NAND2_X1 _12415_ ( .A1(_08957_ ), .A2(_08967_ ), .ZN(_08968_ ) );
NAND2_X1 _12416_ ( .A1(_08963_ ), .A2(_08966_ ), .ZN(_08969_ ) );
AOI21_X4 _12417_ ( .A(_08943_ ), .B1(_08968_ ), .B2(_08969_ ), .ZN(_08970_ ) );
AND3_X1 _12418_ ( .A1(_08941_ ), .A2(_08650_ ), .A3(_08935_ ), .ZN(_08971_ ) );
NOR2_X4 _12419_ ( .A1(_08970_ ), .A2(_08971_ ), .ZN(_08972_ ) );
AND2_X1 _12420_ ( .A1(_08935_ ), .A2(_08604_ ), .ZN(_08973_ ) );
BUF_X4 _12421_ ( .A(_08922_ ), .Z(_08974_ ) );
NAND3_X1 _12422_ ( .A1(_08608_ ), .A2(_08589_ ), .A3(_08974_ ), .ZN(_08975_ ) );
OAI21_X1 _12423_ ( .A(_08975_ ), .B1(dnpc_$_NOT__Y_5_A_$_MUX__Y_A_$_XOR__Y_B ), .B2(_08974_ ), .ZN(_08976_ ) );
XOR2_X1 _12424_ ( .A(_08973_ ), .B(_08976_ ), .Z(_08977_ ) );
INV_X1 _12425_ ( .A(_08977_ ), .ZN(_08978_ ) );
MUX2_X1 _12426_ ( .A(\pc_out[5] ), .B(_08599_ ), .S(_08922_ ), .Z(_08979_ ) );
AND3_X1 _12427_ ( .A1(_08979_ ), .A2(_08595_ ), .A3(_08935_ ), .ZN(_08980_ ) );
AOI21_X1 _12428_ ( .A(_08979_ ), .B1(_08595_ ), .B2(_08935_ ), .ZN(_08981_ ) );
NOR4_X4 _12429_ ( .A1(_08972_ ), .A2(_08978_ ), .A3(_08980_ ), .A4(_08981_ ), .ZN(_08982_ ) );
NOR2_X2 _12430_ ( .A1(_08980_ ), .A2(_08981_ ), .ZN(_08983_ ) );
AND2_X1 _12431_ ( .A1(_08973_ ), .A2(_08976_ ), .ZN(_08984_ ) );
AOI21_X1 _12432_ ( .A(_08980_ ), .B1(_08983_ ), .B2(_08984_ ), .ZN(_08985_ ) );
INV_X1 _12433_ ( .A(_08985_ ), .ZN(_08986_ ) );
OAI21_X2 _12434_ ( .A(_08937_ ), .B1(_08982_ ), .B2(_08986_ ), .ZN(_08987_ ) );
NAND2_X1 _12435_ ( .A1(_08933_ ), .A2(_08936_ ), .ZN(_08988_ ) );
NAND2_X1 _12436_ ( .A1(_08987_ ), .A2(_08988_ ), .ZN(_08989_ ) );
MUX2_X1 _12437_ ( .A(\pc_out[7] ), .B(_08590_ ), .S(_08974_ ), .Z(_08990_ ) );
AND2_X1 _12438_ ( .A1(_08935_ ), .A2(_08582_ ), .ZN(_08991_ ) );
XOR2_X1 _12439_ ( .A(_08990_ ), .B(_08991_ ), .Z(_08992_ ) );
XOR2_X2 _12440_ ( .A(_08989_ ), .B(_08992_ ), .Z(_08993_ ) );
INV_X4 _12441_ ( .A(_08993_ ), .ZN(_08994_ ) );
BUF_X4 _12442_ ( .A(_08994_ ), .Z(_08995_ ) );
BUF_X4 _12443_ ( .A(_08974_ ), .Z(_08996_ ) );
BUF_X4 _12444_ ( .A(_08996_ ), .Z(_08997_ ) );
OAI21_X1 _12445_ ( .A(_08931_ ), .B1(_08995_ ), .B2(_08997_ ), .ZN(_08998_ ) );
AND3_X1 _12446_ ( .A1(\pc_out[3] ), .A2(\pc_out[5] ), .A3(\pc_out[2] ), .ZN(_08999_ ) );
AND2_X2 _12447_ ( .A1(_08999_ ), .A2(\pc_out[4] ), .ZN(_09000_ ) );
NAND2_X1 _12448_ ( .A1(_09000_ ), .A2(_08932_ ), .ZN(_09001_ ) );
INV_X1 _12449_ ( .A(\pc_out[7] ), .ZN(_09002_ ) );
XNOR2_X1 _12450_ ( .A(_09001_ ), .B(_09002_ ), .ZN(_09003_ ) );
NAND3_X1 _12451_ ( .A1(_08906_ ), .A2(_08929_ ), .A3(_09003_ ), .ZN(_09004_ ) );
NAND2_X1 _12452_ ( .A1(_08998_ ), .A2(_09004_ ), .ZN(_09005_ ) );
NAND4_X1 _12453_ ( .A1(_08992_ ), .A2(_08983_ ), .A3(_08937_ ), .A4(_08977_ ), .ZN(_09006_ ) );
NOR2_X1 _12454_ ( .A1(_08972_ ), .A2(_09006_ ), .ZN(_09007_ ) );
AND3_X1 _12455_ ( .A1(_08986_ ), .A2(_08992_ ), .A3(_08937_ ), .ZN(_09008_ ) );
AND2_X1 _12456_ ( .A1(_08990_ ), .A2(_08991_ ), .ZN(_09009_ ) );
AND3_X1 _12457_ ( .A1(_08992_ ), .A2(_08936_ ), .A3(_08933_ ), .ZN(_09010_ ) );
OR3_X4 _12458_ ( .A1(_09008_ ), .A2(_09009_ ), .A3(_09010_ ), .ZN(_09011_ ) );
OR2_X1 _12459_ ( .A1(_09007_ ), .A2(_09011_ ), .ZN(_09012_ ) );
CLKBUF_X2 _12460_ ( .A(_08935_ ), .Z(_09013_ ) );
AND2_X1 _12461_ ( .A1(_09013_ ), .A2(_08678_ ), .ZN(_09014_ ) );
NAND3_X1 _12462_ ( .A1(_08905_ ), .A2(\ifu_rdata[0] ), .A3(\pc_out[8] ), .ZN(_09015_ ) );
OAI21_X1 _12463_ ( .A(_09015_ ), .B1(_08682_ ), .B2(_08921_ ), .ZN(_09016_ ) );
XOR2_X1 _12464_ ( .A(_09014_ ), .B(_09016_ ), .Z(_09017_ ) );
XOR2_X2 _12465_ ( .A(_09012_ ), .B(_09017_ ), .Z(_09018_ ) );
INV_X1 _12466_ ( .A(_09018_ ), .ZN(_09019_ ) );
BUF_X4 _12467_ ( .A(_09019_ ), .Z(_09020_ ) );
OAI21_X1 _12468_ ( .A(_08931_ ), .B1(_09020_ ), .B2(_08997_ ), .ZN(_09021_ ) );
AND3_X1 _12469_ ( .A1(_09000_ ), .A2(\pc_out[7] ), .A3(\pc_out[6] ), .ZN(_09022_ ) );
XNOR2_X1 _12470_ ( .A(_09022_ ), .B(dnpc_$_NOT__Y_1_A_$_MUX__Y_A_$_XOR__Y_B ), .ZN(_09023_ ) );
OR2_X1 _12471_ ( .A1(_08931_ ), .A2(_09023_ ), .ZN(_09024_ ) );
NAND2_X1 _12472_ ( .A1(_09021_ ), .A2(_09024_ ), .ZN(_09025_ ) );
AOI21_X1 _12473_ ( .A(_08575_ ), .B1(_09005_ ), .B2(_09025_ ), .ZN(_09026_ ) );
NAND2_X1 _12474_ ( .A1(_09012_ ), .A2(_09017_ ), .ZN(_09027_ ) );
NAND2_X1 _12475_ ( .A1(_09014_ ), .A2(_09016_ ), .ZN(_09028_ ) );
NAND2_X1 _12476_ ( .A1(_09027_ ), .A2(_09028_ ), .ZN(_09029_ ) );
AND3_X1 _12477_ ( .A1(_08935_ ), .A2(_08636_ ), .A3(_08686_ ), .ZN(_09030_ ) );
NAND3_X1 _12478_ ( .A1(_08905_ ), .A2(\ifu_rdata[0] ), .A3(\pc_out[9] ), .ZN(_09031_ ) );
OAI21_X1 _12479_ ( .A(_09031_ ), .B1(_08692_ ), .B2(_08921_ ), .ZN(_09032_ ) );
XOR2_X1 _12480_ ( .A(_09030_ ), .B(_09032_ ), .Z(_09033_ ) );
XOR2_X1 _12481_ ( .A(_09029_ ), .B(_09033_ ), .Z(_09034_ ) );
BUF_X4 _12482_ ( .A(_09034_ ), .Z(_09035_ ) );
NAND2_X2 _12483_ ( .A1(_08906_ ), .A2(_08928_ ), .ZN(_09036_ ) );
NAND2_X1 _12484_ ( .A1(_09035_ ), .A2(_09036_ ), .ZN(_09037_ ) );
NAND3_X1 _12485_ ( .A1(_09000_ ), .A2(\pc_out[7] ), .A3(\pc_out[6] ), .ZN(_09038_ ) );
NOR2_X1 _12486_ ( .A1(_09038_ ), .A2(dnpc_$_NOT__Y_1_A_$_MUX__Y_A_$_XOR__Y_B ), .ZN(_09039_ ) );
XNOR2_X1 _12487_ ( .A(_09039_ ), .B(\pc_out[9] ), .ZN(_09040_ ) );
OR2_X1 _12488_ ( .A1(_08931_ ), .A2(_09040_ ), .ZN(_09041_ ) );
AOI21_X1 _12489_ ( .A(_08575_ ), .B1(_09037_ ), .B2(_09041_ ), .ZN(_09042_ ) );
NOR2_X1 _12490_ ( .A1(_08982_ ), .A2(_08986_ ), .ZN(_09043_ ) );
XNOR2_X1 _12491_ ( .A(_09043_ ), .B(_08937_ ), .ZN(_09044_ ) );
BUF_X4 _12492_ ( .A(_09044_ ), .Z(_09045_ ) );
BUF_X4 _12493_ ( .A(_09045_ ), .Z(_09046_ ) );
NAND2_X1 _12494_ ( .A1(_09046_ ), .A2(_09036_ ), .ZN(_09047_ ) );
XNOR2_X1 _12495_ ( .A(_09000_ ), .B(dnpc_$_NOT__Y_3_A_$_MUX__Y_A_$_XOR__Y_B ), .ZN(_09048_ ) );
NAND3_X1 _12496_ ( .A1(_08906_ ), .A2(_08929_ ), .A3(_09048_ ), .ZN(_09049_ ) );
AND2_X1 _12497_ ( .A1(_09047_ ), .A2(_09049_ ), .ZN(_09050_ ) );
NOR2_X1 _12498_ ( .A1(_08972_ ), .A2(_08978_ ), .ZN(_09051_ ) );
OR2_X1 _12499_ ( .A1(_09051_ ), .A2(_08984_ ), .ZN(_09052_ ) );
XNOR2_X2 _12500_ ( .A(_09052_ ), .B(_08983_ ), .ZN(_09053_ ) );
BUF_X4 _12501_ ( .A(_09053_ ), .Z(_09054_ ) );
BUF_X4 _12502_ ( .A(_09054_ ), .Z(_09055_ ) );
BUF_X4 _12503_ ( .A(_09055_ ), .Z(_09056_ ) );
OAI21_X1 _12504_ ( .A(_08931_ ), .B1(_09056_ ), .B2(_08997_ ), .ZN(_09057_ ) );
AND2_X1 _12505_ ( .A1(\pc_out[3] ), .A2(\pc_out[2] ), .ZN(_09058_ ) );
INV_X1 _12506_ ( .A(_09058_ ), .ZN(_09059_ ) );
NOR2_X1 _12507_ ( .A1(_09059_ ), .A2(dnpc_$_NOT__Y_5_A_$_MUX__Y_A_$_XOR__Y_B ), .ZN(_09060_ ) );
XNOR2_X1 _12508_ ( .A(_09060_ ), .B(\pc_out[5] ), .ZN(_09061_ ) );
NAND3_X1 _12509_ ( .A1(_08906_ ), .A2(_08929_ ), .A3(_09061_ ), .ZN(_09062_ ) );
NAND2_X1 _12510_ ( .A1(_09057_ ), .A2(_09062_ ), .ZN(_09063_ ) );
AOI21_X1 _12511_ ( .A(_08575_ ), .B1(_09050_ ), .B2(_09063_ ), .ZN(_09064_ ) );
AND3_X1 _12512_ ( .A1(_08968_ ), .A2(_08969_ ), .A3(_08943_ ), .ZN(_09065_ ) );
NOR2_X4 _12513_ ( .A1(_09065_ ), .A2(_08970_ ), .ZN(_09066_ ) );
BUF_X4 _12514_ ( .A(_09066_ ), .Z(_09067_ ) );
BUF_X4 _12515_ ( .A(_09067_ ), .Z(_09068_ ) );
BUF_X4 _12516_ ( .A(_09068_ ), .Z(_09069_ ) );
BUF_X8 _12517_ ( .A(_09069_ ), .Z(_09070_ ) );
BUF_X4 _12518_ ( .A(_09070_ ), .Z(_09071_ ) );
BUF_X2 _12519_ ( .A(_09071_ ), .Z(\alu_result_out[3] ) );
NAND2_X1 _12520_ ( .A1(_09036_ ), .A2(\alu_result_out[3] ), .ZN(_09072_ ) );
XOR2_X1 _12521_ ( .A(\pc_out[3] ), .B(\pc_out[2] ), .Z(_09073_ ) );
INV_X1 _12522_ ( .A(_09073_ ), .ZN(_09074_ ) );
OAI21_X1 _12523_ ( .A(_09072_ ), .B1(_08931_ ), .B2(_09074_ ), .ZN(_09075_ ) );
AND2_X1 _12524_ ( .A1(_09075_ ), .A2(dnpc_$_NOT__Y_A_$_ANDNOT__B_A ), .ZN(_09076_ ) );
INV_X1 _12525_ ( .A(_09076_ ), .ZN(_09077_ ) );
XOR2_X1 _12526_ ( .A(_09058_ ), .B(dnpc_$_NOT__Y_5_A_$_MUX__Y_A_$_XOR__Y_B ), .Z(_09078_ ) );
AOI21_X1 _12527_ ( .A(\u_ifu.reset_sync ), .B1(_08930_ ), .B2(_09078_ ), .ZN(_09079_ ) );
INV_X1 _12528_ ( .A(_09079_ ), .ZN(_09080_ ) );
XNOR2_X1 _12529_ ( .A(_08972_ ), .B(_08977_ ), .ZN(_09081_ ) );
BUF_X4 _12530_ ( .A(_09081_ ), .Z(_09082_ ) );
BUF_X4 _12531_ ( .A(_09082_ ), .Z(_09083_ ) );
BUF_X4 _12532_ ( .A(_09083_ ), .Z(_09084_ ) );
BUF_X4 _12533_ ( .A(_09084_ ), .Z(_09085_ ) );
BUF_X2 _12534_ ( .A(_09085_ ), .Z(\alu_result_out[4] ) );
AOI21_X1 _12535_ ( .A(_08930_ ), .B1(\alu_result_out[4] ), .B2(_08921_ ), .ZN(_09086_ ) );
NOR2_X1 _12536_ ( .A1(_09080_ ), .A2(_09086_ ), .ZN(_00129_ ) );
INV_X1 _12537_ ( .A(_09036_ ), .ZN(_09087_ ) );
XOR2_X1 _12538_ ( .A(_08957_ ), .B(_08967_ ), .Z(_09088_ ) );
BUF_X4 _12539_ ( .A(_09088_ ), .Z(_09089_ ) );
INV_X4 _12540_ ( .A(_09089_ ), .ZN(_09090_ ) );
BUF_X4 _12541_ ( .A(_09090_ ), .Z(_09091_ ) );
BUF_X4 _12542_ ( .A(_09091_ ), .Z(_09092_ ) );
BUF_X4 _12543_ ( .A(_09092_ ), .Z(_09093_ ) );
BUF_X4 _12544_ ( .A(_09093_ ), .Z(_09094_ ) );
BUF_X4 _12545_ ( .A(_09094_ ), .Z(_09095_ ) );
BUF_X2 _12546_ ( .A(_09095_ ), .Z(_09096_ ) );
OAI22_X1 _12547_ ( .A1(_08931_ ), .A2(_08964_ ), .B1(_09087_ ), .B2(_09096_ ), .ZN(_09097_ ) );
INV_X1 _12548_ ( .A(\u_ifu.reset_sync ), .ZN(_09098_ ) );
NAND2_X1 _12549_ ( .A1(_09097_ ), .A2(_09098_ ), .ZN(_09099_ ) );
NAND3_X1 _12550_ ( .A1(_09077_ ), .A2(_00129_ ), .A3(_09099_ ), .ZN(_09100_ ) );
NOR4_X1 _12551_ ( .A1(_09026_ ), .A2(_09042_ ), .A3(_09064_ ), .A4(_09100_ ), .ZN(_00001_ ) );
AOI211_X1 _12552_ ( .A(_09086_ ), .B(_09080_ ), .C1(_09077_ ), .C2(_09099_ ), .ZN(_09101_ ) );
NOR4_X1 _12553_ ( .A1(_09026_ ), .A2(_09042_ ), .A3(_09064_ ), .A4(_09101_ ), .ZN(_00002_ ) );
OR2_X1 _12554_ ( .A1(_09026_ ), .A2(_09064_ ), .ZN(_09102_ ) );
OR2_X1 _12555_ ( .A1(_09102_ ), .A2(_09042_ ), .ZN(_09103_ ) );
NOR3_X1 _12556_ ( .A1(_09103_ ), .A2(_00129_ ), .A3(_09077_ ), .ZN(_00104_ ) );
OR2_X1 _12557_ ( .A1(_00104_ ), .A2(_00001_ ), .ZN(_00003_ ) );
NOR2_X1 _12558_ ( .A1(_09103_ ), .A2(_00129_ ), .ZN(_00004_ ) );
XOR2_X1 _12559_ ( .A(_08951_ ), .B(_08956_ ), .Z(\alu_result_out[1] ) );
INV_X1 _12560_ ( .A(\alu_result_out[1] ), .ZN(_09104_ ) );
BUF_X4 _12561_ ( .A(_08928_ ), .Z(_09105_ ) );
AOI211_X1 _12562_ ( .A(\u_ifu.reset_sync ), .B(_09104_ ), .C1(_08906_ ), .C2(_09105_ ), .ZN(_00101_ ) );
NOR4_X1 _12563_ ( .A1(_09103_ ), .A2(_00129_ ), .A3(_09077_ ), .A4(_09099_ ), .ZN(_00102_ ) );
INV_X1 _12564_ ( .A(_09099_ ), .ZN(_00131_ ) );
NOR4_X1 _12565_ ( .A1(_09102_ ), .A2(_00129_ ), .A3(_00131_ ), .A4(_09042_ ), .ZN(_00107_ ) );
AND2_X1 _12566_ ( .A1(_00107_ ), .A2(_09076_ ), .ZN(_00103_ ) );
NOR4_X1 _12567_ ( .A1(_09102_ ), .A2(_00129_ ), .A3(_09099_ ), .A4(_09042_ ), .ZN(_00105_ ) );
OAI21_X1 _12568_ ( .A(_00004_ ), .B1(_09077_ ), .B2(_09099_ ), .ZN(_09106_ ) );
AOI21_X1 _12569_ ( .A(_09106_ ), .B1(_09077_ ), .B2(_09099_ ), .ZN(_00106_ ) );
BUF_X2 _12570_ ( .A(_09036_ ), .Z(_09107_ ) );
AND3_X1 _12571_ ( .A1(_09107_ ), .A2(_09098_ ), .A3(\pc_out[0] ), .ZN(_00108_ ) );
INV_X1 _12572_ ( .A(fanout_net_8 ), .ZN(_09108_ ) );
BUF_X4 _12573_ ( .A(_09108_ ), .Z(_09109_ ) );
BUF_X4 _12574_ ( .A(_09109_ ), .Z(_09110_ ) );
NOR2_X4 _12575_ ( .A1(_09066_ ), .A2(_09088_ ), .ZN(_09111_ ) );
INV_X1 _12576_ ( .A(_09111_ ), .ZN(_09112_ ) );
NOR2_X1 _12577_ ( .A1(_09081_ ), .A2(_09112_ ), .ZN(_09113_ ) );
AND2_X2 _12578_ ( .A1(_09053_ ), .A2(_09113_ ), .ZN(_09114_ ) );
INV_X1 _12579_ ( .A(_09044_ ), .ZN(_09115_ ) );
AND2_X4 _12580_ ( .A1(_09114_ ), .A2(_09115_ ), .ZN(_09116_ ) );
XNOR2_X2 _12581_ ( .A(_09116_ ), .B(_08995_ ), .ZN(_09117_ ) );
BUF_X4 _12582_ ( .A(_09117_ ), .Z(_09118_ ) );
BUF_X4 _12583_ ( .A(_09083_ ), .Z(_09119_ ) );
NOR2_X4 _12584_ ( .A1(_09066_ ), .A2(_09090_ ), .ZN(_09120_ ) );
BUF_X4 _12585_ ( .A(_09120_ ), .Z(_09121_ ) );
BUF_X8 _12586_ ( .A(_09121_ ), .Z(_09122_ ) );
BUF_X8 _12587_ ( .A(_09122_ ), .Z(_09123_ ) );
INV_X4 _12588_ ( .A(_09123_ ), .ZN(_09124_ ) );
NOR2_X4 _12589_ ( .A1(_09119_ ), .A2(_09124_ ), .ZN(_09125_ ) );
INV_X1 _12590_ ( .A(_09125_ ), .ZN(_09126_ ) );
NOR2_X4 _12591_ ( .A1(_09055_ ), .A2(_09126_ ), .ZN(_09127_ ) );
INV_X1 _12592_ ( .A(_09127_ ), .ZN(_09128_ ) );
XNOR2_X2 _12593_ ( .A(_09114_ ), .B(_09045_ ), .ZN(_09129_ ) );
INV_X1 _12594_ ( .A(_09129_ ), .ZN(_09130_ ) );
NOR3_X2 _12595_ ( .A1(_09118_ ), .A2(_09128_ ), .A3(_09130_ ), .ZN(_09131_ ) );
INV_X1 _12596_ ( .A(_09131_ ), .ZN(_09132_ ) );
AND2_X4 _12597_ ( .A1(_09116_ ), .A2(_08994_ ), .ZN(_09133_ ) );
XNOR2_X2 _12598_ ( .A(_09133_ ), .B(_09019_ ), .ZN(_09134_ ) );
BUF_X4 _12599_ ( .A(_09134_ ), .Z(_09135_ ) );
NOR2_X4 _12600_ ( .A1(_09132_ ), .A2(_09135_ ), .ZN(_09136_ ) );
AND2_X4 _12601_ ( .A1(_09133_ ), .A2(_09019_ ), .ZN(_09137_ ) );
INV_X2 _12602_ ( .A(_09034_ ), .ZN(_09138_ ) );
XNOR2_X1 _12603_ ( .A(_09137_ ), .B(_09138_ ), .ZN(_09139_ ) );
BUF_X8 _12604_ ( .A(_09139_ ), .Z(_09140_ ) );
BUF_X4 _12605_ ( .A(_09140_ ), .Z(_09141_ ) );
AND2_X1 _12606_ ( .A1(_09136_ ), .A2(_09141_ ), .ZN(_09142_ ) );
OAI21_X1 _12607_ ( .A(_09110_ ), .B1(_09142_ ), .B2(\u_lsu.pmem[4388] ), .ZN(_09143_ ) );
AND2_X4 _12608_ ( .A1(_09137_ ), .A2(_09138_ ), .ZN(_09144_ ) );
BUF_X4 _12609_ ( .A(_09144_ ), .Z(_09145_ ) );
INV_X1 _12610_ ( .A(_08605_ ), .ZN(_09146_ ) );
NOR2_X4 _12611_ ( .A1(_09145_ ), .A2(_09146_ ), .ZN(_09147_ ) );
BUF_X4 _12612_ ( .A(_09147_ ), .Z(_09148_ ) );
INV_X1 _12613_ ( .A(_09148_ ), .ZN(_09149_ ) );
AOI21_X1 _12614_ ( .A(_09143_ ), .B1(_09142_ ), .B2(_09149_ ), .ZN(_00109_ ) );
MUX2_X1 _12615_ ( .A(\pc_out[19] ), .B(_08752_ ), .S(_08996_ ), .Z(_09150_ ) );
AND2_X1 _12616_ ( .A1(_09013_ ), .A2(_08748_ ), .ZN(_09151_ ) );
XOR2_X1 _12617_ ( .A(_09150_ ), .B(_09151_ ), .Z(_09152_ ) );
MUX2_X1 _12618_ ( .A(\pc_out[18] ), .B(_08762_ ), .S(_08996_ ), .Z(_09153_ ) );
AND3_X1 _12619_ ( .A1(_09013_ ), .A2(_08637_ ), .A3(_08756_ ), .ZN(_09154_ ) );
XOR2_X1 _12620_ ( .A(_09153_ ), .B(_09154_ ), .Z(_09155_ ) );
AND2_X1 _12621_ ( .A1(_09152_ ), .A2(_09155_ ), .ZN(_09156_ ) );
AND2_X1 _12622_ ( .A1(_08779_ ), .A2(_08589_ ), .ZN(_09157_ ) );
MUX2_X1 _12623_ ( .A(\pc_out[17] ), .B(_09157_ ), .S(_08974_ ), .Z(_09158_ ) );
AND3_X1 _12624_ ( .A1(_09013_ ), .A2(_08636_ ), .A3(_08776_ ), .ZN(_09159_ ) );
XOR2_X1 _12625_ ( .A(_09158_ ), .B(_09159_ ), .Z(_09160_ ) );
AND3_X1 _12626_ ( .A1(_08921_ ), .A2(_08959_ ), .A3(\ifu_rdata[2] ), .ZN(_09161_ ) );
AOI21_X1 _12627_ ( .A(_09161_ ), .B1(_09013_ ), .B2(_08768_ ), .ZN(_09162_ ) );
NAND3_X1 _12628_ ( .A1(_08905_ ), .A2(\ifu_rdata[0] ), .A3(dnpc_$_MUX__Y_15_A_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_09163_ ) );
OAI21_X1 _12629_ ( .A(_09163_ ), .B1(_08772_ ), .B2(_08921_ ), .ZN(_09164_ ) );
NOR2_X1 _12630_ ( .A1(_09162_ ), .A2(_09164_ ), .ZN(_09165_ ) );
AND2_X1 _12631_ ( .A1(_09160_ ), .A2(_09165_ ), .ZN(_09166_ ) );
AOI21_X1 _12632_ ( .A(_09166_ ), .B1(_09159_ ), .B2(_09158_ ), .ZN(_09167_ ) );
INV_X1 _12633_ ( .A(_09167_ ), .ZN(_09168_ ) );
AND2_X1 _12634_ ( .A1(_09156_ ), .A2(_09168_ ), .ZN(_09169_ ) );
AND2_X1 _12635_ ( .A1(_09150_ ), .A2(_09151_ ), .ZN(_09170_ ) );
AND2_X1 _12636_ ( .A1(_09153_ ), .A2(_09154_ ), .ZN(_09171_ ) );
AND2_X1 _12637_ ( .A1(_09152_ ), .A2(_09171_ ), .ZN(_09172_ ) );
NOR3_X1 _12638_ ( .A1(_09169_ ), .A2(_09170_ ), .A3(_09172_ ), .ZN(_09173_ ) );
MUX2_X1 _12639_ ( .A(\pc_out[23] ), .B(_08808_ ), .S(_08996_ ), .Z(_09174_ ) );
CLKBUF_X2 _12640_ ( .A(_09013_ ), .Z(_09175_ ) );
AND2_X1 _12641_ ( .A1(_09175_ ), .A2(_08804_ ), .ZN(_09176_ ) );
XNOR2_X1 _12642_ ( .A(_09174_ ), .B(_09176_ ), .ZN(_09177_ ) );
AND3_X1 _12643_ ( .A1(_08905_ ), .A2(\ifu_rdata[0] ), .A3(\pc_out[22] ), .ZN(_09178_ ) );
AOI21_X1 _12644_ ( .A(_09178_ ), .B1(_08813_ ), .B2(_08996_ ), .ZN(_09179_ ) );
NAND3_X1 _12645_ ( .A1(_08944_ ), .A2(_08818_ ), .A3(_08934_ ), .ZN(_09180_ ) );
XNOR2_X1 _12646_ ( .A(_09179_ ), .B(_09180_ ), .ZN(_09181_ ) );
NOR2_X1 _12647_ ( .A1(_09177_ ), .A2(_09181_ ), .ZN(_09182_ ) );
INV_X1 _12648_ ( .A(_09182_ ), .ZN(_09183_ ) );
MUX2_X1 _12649_ ( .A(\pc_out[21] ), .B(_08799_ ), .S(_08996_ ), .Z(_09184_ ) );
AND2_X1 _12650_ ( .A1(_09013_ ), .A2(_08795_ ), .ZN(_09185_ ) );
XOR2_X1 _12651_ ( .A(_09184_ ), .B(_09185_ ), .Z(_09186_ ) );
INV_X1 _12652_ ( .A(_09186_ ), .ZN(_09187_ ) );
INV_X1 _12653_ ( .A(dnpc_$_MUX__Y_11_A_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_09188_ ) );
MUX2_X1 _12654_ ( .A(_09188_ ), .B(_08786_ ), .S(_08996_ ), .Z(_09189_ ) );
AND3_X1 _12655_ ( .A1(_09175_ ), .A2(_08637_ ), .A3(_08789_ ), .ZN(_09190_ ) );
XNOR2_X1 _12656_ ( .A(_09189_ ), .B(_09190_ ), .ZN(_09191_ ) );
NOR4_X1 _12657_ ( .A1(_09173_ ), .A2(_09183_ ), .A3(_09187_ ), .A4(_09191_ ), .ZN(_09192_ ) );
AND2_X1 _12658_ ( .A1(_09174_ ), .A2(_09176_ ), .ZN(_09193_ ) );
NAND2_X1 _12659_ ( .A1(_09184_ ), .A2(_09185_ ), .ZN(_09194_ ) );
NAND2_X1 _12660_ ( .A1(_09189_ ), .A2(_09190_ ), .ZN(_09195_ ) );
OAI21_X1 _12661_ ( .A(_09194_ ), .B1(_09187_ ), .B2(_09195_ ), .ZN(_09196_ ) );
AND2_X1 _12662_ ( .A1(_09196_ ), .A2(_09182_ ), .ZN(_09197_ ) );
NOR3_X1 _12663_ ( .A1(_09177_ ), .A2(_09180_ ), .A3(_09179_ ), .ZN(_09198_ ) );
NOR4_X1 _12664_ ( .A1(_09192_ ), .A2(_09193_ ), .A3(_09197_ ), .A4(_09198_ ), .ZN(_09199_ ) );
MUX2_X1 _12665_ ( .A(\pc_out[15] ), .B(_08723_ ), .S(_08996_ ), .Z(_09200_ ) );
NAND4_X1 _12666_ ( .A1(_08944_ ), .A2(_08718_ ), .A3(_08636_ ), .A4(_08934_ ), .ZN(_09201_ ) );
OAI21_X1 _12667_ ( .A(_09201_ ), .B1(_08587_ ), .B2(_08909_ ), .ZN(_09202_ ) );
NAND2_X1 _12668_ ( .A1(_09200_ ), .A2(_09202_ ), .ZN(_09203_ ) );
AND2_X1 _12669_ ( .A1(_09013_ ), .A2(_08741_ ), .ZN(_09204_ ) );
MUX2_X1 _12670_ ( .A(\pc_out[14] ), .B(_08737_ ), .S(_08974_ ), .Z(_09205_ ) );
OAI211_X1 _12671_ ( .A(_09204_ ), .B(_09205_ ), .C1(_09200_ ), .C2(_09202_ ), .ZN(_09206_ ) );
MUX2_X1 _12672_ ( .A(\pc_out[11] ), .B(_08669_ ), .S(_08974_ ), .Z(_09207_ ) );
NAND4_X1 _12673_ ( .A1(_08905_ ), .A2(_08924_ ), .A3(\ifu_rdata[2] ), .A4(\ifu_rdata[0] ), .ZN(_09208_ ) );
NAND3_X1 _12674_ ( .A1(_08905_ ), .A2(\ifu_rdata[7] ), .A3(_08902_ ), .ZN(_09209_ ) );
AND2_X1 _12675_ ( .A1(_09208_ ), .A2(_09209_ ), .ZN(_09210_ ) );
OAI21_X1 _12676_ ( .A(_09210_ ), .B1(_08953_ ), .B2(_08673_ ), .ZN(_09211_ ) );
XNOR2_X1 _12677_ ( .A(_09207_ ), .B(_09211_ ), .ZN(_09212_ ) );
MUX2_X1 _12678_ ( .A(\pc_out[10] ), .B(_08697_ ), .S(_08974_ ), .Z(_09213_ ) );
AND3_X1 _12679_ ( .A1(_08944_ ), .A2(_08704_ ), .A3(_08934_ ), .ZN(_09214_ ) );
XNOR2_X1 _12680_ ( .A(_09213_ ), .B(_09214_ ), .ZN(_09215_ ) );
NAND3_X1 _12681_ ( .A1(_09033_ ), .A2(_09014_ ), .A3(_09016_ ), .ZN(_09216_ ) );
NAND2_X1 _12682_ ( .A1(_09030_ ), .A2(_09032_ ), .ZN(_09217_ ) );
AOI211_X1 _12683_ ( .A(_09212_ ), .B(_09215_ ), .C1(_09216_ ), .C2(_09217_ ), .ZN(_09218_ ) );
AND2_X1 _12684_ ( .A1(_09207_ ), .A2(_09211_ ), .ZN(_09219_ ) );
AND2_X1 _12685_ ( .A1(_09213_ ), .A2(_09214_ ), .ZN(_09220_ ) );
INV_X1 _12686_ ( .A(_09220_ ), .ZN(_09221_ ) );
NOR2_X1 _12687_ ( .A1(_09212_ ), .A2(_09221_ ), .ZN(_09222_ ) );
NOR3_X1 _12688_ ( .A1(_09218_ ), .A2(_09219_ ), .A3(_09222_ ), .ZN(_09223_ ) );
XNOR2_X1 _12689_ ( .A(_09200_ ), .B(_09202_ ), .ZN(_09224_ ) );
XNOR2_X1 _12690_ ( .A(_09205_ ), .B(_09204_ ), .ZN(_09225_ ) );
NOR2_X1 _12691_ ( .A1(_09224_ ), .A2(_09225_ ), .ZN(_09226_ ) );
MUX2_X1 _12692_ ( .A(\pc_out[12] ), .B(_08728_ ), .S(_08974_ ), .Z(_09227_ ) );
AND2_X1 _12693_ ( .A1(_09013_ ), .A2(_08732_ ), .ZN(_09228_ ) );
XNOR2_X1 _12694_ ( .A(_09227_ ), .B(_09228_ ), .ZN(_09229_ ) );
MUX2_X1 _12695_ ( .A(\pc_out[13] ), .B(_08714_ ), .S(_08974_ ), .Z(_09230_ ) );
AND2_X1 _12696_ ( .A1(_09013_ ), .A2(_08710_ ), .ZN(_09231_ ) );
XNOR2_X1 _12697_ ( .A(_09230_ ), .B(_09231_ ), .ZN(_09232_ ) );
NOR2_X1 _12698_ ( .A1(_09229_ ), .A2(_09232_ ), .ZN(_09233_ ) );
AND2_X1 _12699_ ( .A1(_09226_ ), .A2(_09233_ ), .ZN(_09234_ ) );
INV_X1 _12700_ ( .A(_09234_ ), .ZN(_09235_ ) );
OAI211_X1 _12701_ ( .A(_09203_ ), .B(_09206_ ), .C1(_09223_ ), .C2(_09235_ ), .ZN(_09236_ ) );
OAI211_X1 _12702_ ( .A(_09228_ ), .B(_09227_ ), .C1(_09230_ ), .C2(_09231_ ), .ZN(_09237_ ) );
NAND2_X1 _12703_ ( .A1(_09230_ ), .A2(_09231_ ), .ZN(_09238_ ) );
NAND2_X1 _12704_ ( .A1(_09237_ ), .A2(_09238_ ), .ZN(_09239_ ) );
AOI21_X1 _12705_ ( .A(_09236_ ), .B1(_09226_ ), .B2(_09239_ ), .ZN(_09240_ ) );
NAND2_X1 _12706_ ( .A1(_09033_ ), .A2(_09017_ ), .ZN(_09241_ ) );
NOR3_X1 _12707_ ( .A1(_09241_ ), .A2(_09212_ ), .A3(_09215_ ), .ZN(_09242_ ) );
OAI211_X1 _12708_ ( .A(_09234_ ), .B(_09242_ ), .C1(_09007_ ), .C2(_09011_ ), .ZN(_09243_ ) );
NAND2_X1 _12709_ ( .A1(_09240_ ), .A2(_09243_ ), .ZN(_09244_ ) );
NOR3_X1 _12710_ ( .A1(_09183_ ), .A2(_09187_ ), .A3(_09191_ ), .ZN(_09245_ ) );
XOR2_X1 _12711_ ( .A(_09162_ ), .B(_09164_ ), .Z(_09246_ ) );
AND2_X1 _12712_ ( .A1(_09160_ ), .A2(_09246_ ), .ZN(_09247_ ) );
AND2_X1 _12713_ ( .A1(_09156_ ), .A2(_09247_ ), .ZN(_09248_ ) );
NAND3_X1 _12714_ ( .A1(_09244_ ), .A2(_09245_ ), .A3(_09248_ ), .ZN(_09249_ ) );
NAND2_X1 _12715_ ( .A1(_09199_ ), .A2(_09249_ ), .ZN(_09250_ ) );
MUX2_X1 _12716_ ( .A(\pc_out[27] ), .B(_08881_ ), .S(_08997_ ), .Z(_09251_ ) );
AND3_X1 _12717_ ( .A1(_09175_ ), .A2(_08687_ ), .A3(_08884_ ), .ZN(_09252_ ) );
XOR2_X1 _12718_ ( .A(_09251_ ), .B(_09252_ ), .Z(_09253_ ) );
MUX2_X1 _12719_ ( .A(\pc_out[26] ), .B(_08895_ ), .S(_08997_ ), .Z(_09254_ ) );
AND2_X1 _12720_ ( .A1(_09175_ ), .A2(_08890_ ), .ZN(_09255_ ) );
XOR2_X1 _12721_ ( .A(_09254_ ), .B(_09255_ ), .Z(_09256_ ) );
MUX2_X1 _12722_ ( .A(\pc_out[24] ), .B(_08871_ ), .S(_08996_ ), .Z(_09257_ ) );
AND3_X1 _12723_ ( .A1(_08876_ ), .A2(_08944_ ), .A3(_08934_ ), .ZN(_09258_ ) );
XOR2_X1 _12724_ ( .A(_09257_ ), .B(_09258_ ), .Z(_09259_ ) );
MUX2_X1 _12725_ ( .A(\pc_out[25] ), .B(_08866_ ), .S(_08996_ ), .Z(_09260_ ) );
AND2_X1 _12726_ ( .A1(_09175_ ), .A2(_08862_ ), .ZN(_09261_ ) );
XOR2_X1 _12727_ ( .A(_09260_ ), .B(_09261_ ), .Z(_09262_ ) );
AND2_X1 _12728_ ( .A1(_09259_ ), .A2(_09262_ ), .ZN(_09263_ ) );
NAND4_X1 _12729_ ( .A1(_09250_ ), .A2(_09253_ ), .A3(_09256_ ), .A4(_09263_ ), .ZN(_09264_ ) );
AND2_X1 _12730_ ( .A1(_09254_ ), .A2(_09255_ ), .ZN(_09265_ ) );
AND2_X1 _12731_ ( .A1(_09253_ ), .A2(_09265_ ), .ZN(_09266_ ) );
AND2_X1 _12732_ ( .A1(_09257_ ), .A2(_09258_ ), .ZN(_09267_ ) );
AND2_X1 _12733_ ( .A1(_09262_ ), .A2(_09267_ ), .ZN(_09268_ ) );
AOI21_X1 _12734_ ( .A(_09268_ ), .B1(_09261_ ), .B2(_09260_ ), .ZN(_09269_ ) );
INV_X1 _12735_ ( .A(_09269_ ), .ZN(_09270_ ) );
AND3_X1 _12736_ ( .A1(_09270_ ), .A2(_09253_ ), .A3(_09256_ ), .ZN(_09271_ ) );
AOI211_X1 _12737_ ( .A(_09266_ ), .B(_09271_ ), .C1(_09252_ ), .C2(_09251_ ), .ZN(_09272_ ) );
AND2_X1 _12738_ ( .A1(_09264_ ), .A2(_09272_ ), .ZN(_09273_ ) );
AND2_X1 _12739_ ( .A1(_09175_ ), .A2(_08824_ ), .ZN(_09274_ ) );
NAND3_X1 _12740_ ( .A1(_08905_ ), .A2(\ifu_rdata[0] ), .A3(\pc_out[29] ), .ZN(_09275_ ) );
OAI21_X1 _12741_ ( .A(_09275_ ), .B1(_08828_ ), .B2(_08921_ ), .ZN(_09276_ ) );
XNOR2_X1 _12742_ ( .A(_09274_ ), .B(_09276_ ), .ZN(_09277_ ) );
MUX2_X1 _12743_ ( .A(\pc_out[28] ), .B(_08842_ ), .S(_08997_ ), .Z(_09278_ ) );
AND2_X1 _12744_ ( .A1(_09175_ ), .A2(_08846_ ), .ZN(_09279_ ) );
XNOR2_X1 _12745_ ( .A(_09278_ ), .B(_09279_ ), .ZN(_09280_ ) );
OR3_X1 _12746_ ( .A1(_09273_ ), .A2(_09277_ ), .A3(_09280_ ), .ZN(_09281_ ) );
NAND3_X1 _12747_ ( .A1(_09276_ ), .A2(_08824_ ), .A3(_09175_ ), .ZN(_09282_ ) );
OAI211_X1 _12748_ ( .A(_09278_ ), .B(_09279_ ), .C1(_09274_ ), .C2(_09276_ ), .ZN(_09283_ ) );
AND3_X1 _12749_ ( .A1(_09281_ ), .A2(_09282_ ), .A3(_09283_ ), .ZN(_09284_ ) );
AND2_X1 _12750_ ( .A1(_09175_ ), .A2(_08856_ ), .ZN(_09285_ ) );
NAND3_X1 _12751_ ( .A1(_08850_ ), .A2(_08611_ ), .A3(_08997_ ), .ZN(_09286_ ) );
NAND3_X1 _12752_ ( .A1(_08905_ ), .A2(\ifu_rdata[0] ), .A3(\pc_out[30] ), .ZN(_09287_ ) );
NAND2_X1 _12753_ ( .A1(_09286_ ), .A2(_09287_ ), .ZN(_09288_ ) );
XNOR2_X1 _12754_ ( .A(_09285_ ), .B(_09288_ ), .ZN(_09289_ ) );
XOR2_X1 _12755_ ( .A(_09284_ ), .B(_09289_ ), .Z(\alu_result_out[30] ) );
BUF_X4 _12756_ ( .A(_09036_ ), .Z(_09290_ ) );
BUF_X4 _12757_ ( .A(_08930_ ), .Z(_09291_ ) );
AND2_X1 _12758_ ( .A1(\pc_out[11] ), .A2(\pc_out[10] ), .ZN(_09292_ ) );
AND3_X1 _12759_ ( .A1(_09292_ ), .A2(\pc_out[13] ), .A3(\pc_out[12] ), .ZN(_09293_ ) );
AND2_X1 _12760_ ( .A1(\pc_out[15] ), .A2(\pc_out[14] ), .ZN(_09294_ ) );
AND4_X1 _12761_ ( .A1(\pc_out[17] ), .A2(_09293_ ), .A3(\pc_out[16] ), .A4(_09294_ ), .ZN(_09295_ ) );
AND4_X1 _12762_ ( .A1(\pc_out[7] ), .A2(\pc_out[6] ), .A3(\pc_out[9] ), .A4(\pc_out[8] ), .ZN(_09296_ ) );
AND2_X2 _12763_ ( .A1(_09000_ ), .A2(_09296_ ), .ZN(_09297_ ) );
AND2_X1 _12764_ ( .A1(_09295_ ), .A2(_09297_ ), .ZN(_09298_ ) );
AND2_X1 _12765_ ( .A1(\pc_out[19] ), .A2(\pc_out[18] ), .ZN(_09299_ ) );
AND3_X1 _12766_ ( .A1(_09299_ ), .A2(\pc_out[21] ), .A3(\pc_out[20] ), .ZN(_09300_ ) );
AND2_X1 _12767_ ( .A1(\pc_out[23] ), .A2(\pc_out[22] ), .ZN(_09301_ ) );
AND4_X1 _12768_ ( .A1(\pc_out[25] ), .A2(_09300_ ), .A3(\pc_out[24] ), .A4(_09301_ ), .ZN(_09302_ ) );
AND4_X1 _12769_ ( .A1(\pc_out[29] ), .A2(\pc_out[28] ), .A3(\pc_out[27] ), .A4(\pc_out[26] ), .ZN(_09303_ ) );
AND3_X1 _12770_ ( .A1(_09298_ ), .A2(_09302_ ), .A3(_09303_ ), .ZN(_09304_ ) );
XNOR2_X1 _12771_ ( .A(_09304_ ), .B(dnpc_$_MUX__Y_1_A_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_09305_ ) );
AOI22_X1 _12772_ ( .A1(\alu_result_out[30] ), .A2(_09290_ ), .B1(_09291_ ), .B2(_09305_ ), .ZN(_09306_ ) );
NOR2_X1 _12773_ ( .A1(_09306_ ), .A2(\u_ifu.reset_sync ), .ZN(_00110_ ) );
AOI21_X1 _12774_ ( .A(_09280_ ), .B1(_09264_ ), .B2(_09272_ ), .ZN(_09307_ ) );
AND2_X1 _12775_ ( .A1(_09278_ ), .A2(_09279_ ), .ZN(_09308_ ) );
OR2_X1 _12776_ ( .A1(_09307_ ), .A2(_09308_ ), .ZN(_09309_ ) );
XNOR2_X1 _12777_ ( .A(_09309_ ), .B(_09277_ ), .ZN(\alu_result_out[29] ) );
NAND2_X1 _12778_ ( .A1(\alu_result_out[29] ), .A2(_09107_ ), .ZN(_09310_ ) );
BUF_X1 _12779_ ( .A(_08931_ ), .Z(jump_en ) );
AND2_X1 _12780_ ( .A1(_09298_ ), .A2(_09302_ ), .ZN(_09311_ ) );
AND3_X1 _12781_ ( .A1(_09311_ ), .A2(\pc_out[27] ), .A3(\pc_out[26] ), .ZN(_09312_ ) );
INV_X1 _12782_ ( .A(_09312_ ), .ZN(_09313_ ) );
NOR2_X1 _12783_ ( .A1(_09313_ ), .A2(dnpc_$_MUX__Y_3_A_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_09314_ ) );
XNOR2_X1 _12784_ ( .A(_09314_ ), .B(\pc_out[29] ), .ZN(_09315_ ) );
OR2_X1 _12785_ ( .A1(jump_en ), .A2(_09315_ ), .ZN(_09316_ ) );
AOI21_X1 _12786_ ( .A(\u_ifu.reset_sync ), .B1(_09310_ ), .B2(_09316_ ), .ZN(_00111_ ) );
NAND2_X1 _12787_ ( .A1(_09244_ ), .A2(_09248_ ), .ZN(_09317_ ) );
NAND2_X1 _12788_ ( .A1(_09317_ ), .A2(_09173_ ), .ZN(_09318_ ) );
XNOR2_X1 _12789_ ( .A(_09318_ ), .B(_09191_ ), .ZN(\alu_result_out[20] ) );
NAND3_X1 _12790_ ( .A1(_09295_ ), .A2(_09299_ ), .A3(_09297_ ), .ZN(_09319_ ) );
XNOR2_X1 _12791_ ( .A(_09319_ ), .B(_09188_ ), .ZN(_09320_ ) );
AOI22_X1 _12792_ ( .A1(\alu_result_out[20] ), .A2(_09290_ ), .B1(_09291_ ), .B2(_09320_ ), .ZN(_09321_ ) );
NOR2_X1 _12793_ ( .A1(_09321_ ), .A2(\u_ifu.reset_sync ), .ZN(_00112_ ) );
AOI21_X1 _12794_ ( .A(_09168_ ), .B1(_09244_ ), .B2(_09247_ ), .ZN(_09322_ ) );
XNOR2_X1 _12795_ ( .A(_09153_ ), .B(_09154_ ), .ZN(_09323_ ) );
NOR2_X1 _12796_ ( .A1(_09322_ ), .A2(_09323_ ), .ZN(_09324_ ) );
NOR2_X1 _12797_ ( .A1(_09324_ ), .A2(_09171_ ), .ZN(_09325_ ) );
XNOR2_X1 _12798_ ( .A(_09325_ ), .B(_09152_ ), .ZN(\alu_result_out[19] ) );
NAND2_X1 _12799_ ( .A1(\alu_result_out[19] ), .A2(_09107_ ), .ZN(_09326_ ) );
INV_X1 _12800_ ( .A(dnpc_$_MUX__Y_13_A_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_09327_ ) );
AND3_X1 _12801_ ( .A1(_09295_ ), .A2(_09327_ ), .A3(_09297_ ), .ZN(_09328_ ) );
XNOR2_X1 _12802_ ( .A(_09328_ ), .B(\pc_out[19] ), .ZN(_09329_ ) );
OR2_X1 _12803_ ( .A1(jump_en ), .A2(_09329_ ), .ZN(_09330_ ) );
AOI21_X1 _12804_ ( .A(\u_ifu.reset_sync ), .B1(_09326_ ), .B2(_09330_ ), .ZN(_00113_ ) );
XNOR2_X1 _12805_ ( .A(_09322_ ), .B(_09155_ ), .ZN(\alu_result_out[18] ) );
XNOR2_X1 _12806_ ( .A(_09298_ ), .B(dnpc_$_MUX__Y_13_A_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_09331_ ) );
AOI22_X1 _12807_ ( .A1(\alu_result_out[18] ), .A2(_09290_ ), .B1(_09291_ ), .B2(_09331_ ), .ZN(_09332_ ) );
NOR2_X1 _12808_ ( .A1(_09332_ ), .A2(\u_ifu.reset_sync ), .ZN(_00114_ ) );
INV_X1 _12809_ ( .A(_09246_ ), .ZN(_09333_ ) );
OAI211_X1 _12810_ ( .A(_09234_ ), .B(_09242_ ), .C1(_09007_ ), .C2(_09011_ ), .ZN(_09334_ ) );
AOI21_X1 _12811_ ( .A(_09333_ ), .B1(_09240_ ), .B2(_09334_ ), .ZN(_09335_ ) );
NOR2_X1 _12812_ ( .A1(_09335_ ), .A2(_09165_ ), .ZN(_09336_ ) );
XNOR2_X1 _12813_ ( .A(_09336_ ), .B(_09160_ ), .ZN(\alu_result_out[17] ) );
NAND2_X1 _12814_ ( .A1(\alu_result_out[17] ), .A2(_09107_ ), .ZN(_09337_ ) );
NAND3_X1 _12815_ ( .A1(_09297_ ), .A2(_09294_ ), .A3(_09293_ ), .ZN(_09338_ ) );
NOR2_X1 _12816_ ( .A1(_09338_ ), .A2(dnpc_$_MUX__Y_15_A_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_09339_ ) );
XNOR2_X1 _12817_ ( .A(_09339_ ), .B(\pc_out[17] ), .ZN(_09340_ ) );
OR2_X1 _12818_ ( .A1(jump_en ), .A2(_09340_ ), .ZN(_09341_ ) );
AOI21_X1 _12819_ ( .A(\u_ifu.reset_sync ), .B1(_09337_ ), .B2(_09341_ ), .ZN(_00115_ ) );
XNOR2_X1 _12820_ ( .A(_09244_ ), .B(_09333_ ), .ZN(\alu_result_out[16] ) );
AND3_X1 _12821_ ( .A1(_09297_ ), .A2(_09294_ ), .A3(_09293_ ), .ZN(_09342_ ) );
XNOR2_X1 _12822_ ( .A(_09342_ ), .B(dnpc_$_MUX__Y_15_A_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_09343_ ) );
AOI22_X1 _12823_ ( .A1(\alu_result_out[16] ), .A2(_09290_ ), .B1(_09291_ ), .B2(_09343_ ), .ZN(_09344_ ) );
NOR2_X1 _12824_ ( .A1(_09344_ ), .A2(\u_ifu.reset_sync ), .ZN(_00116_ ) );
OAI21_X1 _12825_ ( .A(_09242_ ), .B1(_09007_ ), .B2(_09011_ ), .ZN(_09345_ ) );
AOI211_X1 _12826_ ( .A(_09232_ ), .B(_09229_ ), .C1(_09345_ ), .C2(_09223_ ), .ZN(_09346_ ) );
NOR2_X1 _12827_ ( .A1(_09346_ ), .A2(_09239_ ), .ZN(_09347_ ) );
NOR2_X1 _12828_ ( .A1(_09347_ ), .A2(_09225_ ), .ZN(_09348_ ) );
AND2_X1 _12829_ ( .A1(_09205_ ), .A2(_09204_ ), .ZN(_09349_ ) );
OR2_X1 _12830_ ( .A1(_09348_ ), .A2(_09349_ ), .ZN(_09350_ ) );
XNOR2_X1 _12831_ ( .A(_09350_ ), .B(_09224_ ), .ZN(\alu_result_out[15] ) );
NAND2_X1 _12832_ ( .A1(\alu_result_out[15] ), .A2(_09107_ ), .ZN(_09351_ ) );
INV_X1 _12833_ ( .A(dnpc_$_MUX__Y_17_A_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_09352_ ) );
AND3_X1 _12834_ ( .A1(_09297_ ), .A2(_09352_ ), .A3(_09293_ ), .ZN(_09353_ ) );
XNOR2_X1 _12835_ ( .A(_09353_ ), .B(\pc_out[15] ), .ZN(_09354_ ) );
OR2_X1 _12836_ ( .A1(jump_en ), .A2(_09354_ ), .ZN(_09355_ ) );
AOI21_X1 _12837_ ( .A(\u_ifu.reset_sync ), .B1(_09351_ ), .B2(_09355_ ), .ZN(_00117_ ) );
XOR2_X1 _12838_ ( .A(_09347_ ), .B(_09225_ ), .Z(\alu_result_out[14] ) );
AND2_X1 _12839_ ( .A1(_09297_ ), .A2(_09293_ ), .ZN(_09356_ ) );
XNOR2_X1 _12840_ ( .A(_09356_ ), .B(dnpc_$_MUX__Y_17_A_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_09357_ ) );
AOI22_X1 _12841_ ( .A1(\alu_result_out[14] ), .A2(_09290_ ), .B1(_09291_ ), .B2(_09357_ ), .ZN(_09358_ ) );
NOR2_X1 _12842_ ( .A1(_09358_ ), .A2(\u_ifu.reset_sync ), .ZN(_00118_ ) );
AOI21_X1 _12843_ ( .A(_09229_ ), .B1(_09345_ ), .B2(_09223_ ), .ZN(_09359_ ) );
AND2_X1 _12844_ ( .A1(_09227_ ), .A2(_09228_ ), .ZN(_09360_ ) );
OR2_X1 _12845_ ( .A1(_09359_ ), .A2(_09360_ ), .ZN(_09361_ ) );
XNOR2_X1 _12846_ ( .A(_09361_ ), .B(_09232_ ), .ZN(\alu_result_out[13] ) );
AND3_X1 _12847_ ( .A1(_09022_ ), .A2(\pc_out[9] ), .A3(\pc_out[8] ), .ZN(_09362_ ) );
AND3_X1 _12848_ ( .A1(_09362_ ), .A2(\pc_out[12] ), .A3(_09292_ ), .ZN(_09363_ ) );
XOR2_X1 _12849_ ( .A(_09363_ ), .B(\pc_out[13] ), .Z(_09364_ ) );
AOI22_X1 _12850_ ( .A1(\alu_result_out[13] ), .A2(_09290_ ), .B1(_09291_ ), .B2(_09364_ ), .ZN(_09365_ ) );
NOR2_X1 _12851_ ( .A1(_09365_ ), .A2(\u_ifu.reset_sync ), .ZN(_00119_ ) );
NAND2_X1 _12852_ ( .A1(_09345_ ), .A2(_09223_ ), .ZN(_09366_ ) );
XNOR2_X1 _12853_ ( .A(_09366_ ), .B(_09229_ ), .ZN(\alu_result_out[12] ) );
AND3_X1 _12854_ ( .A1(_09000_ ), .A2(_09292_ ), .A3(_09296_ ), .ZN(_09367_ ) );
XOR2_X1 _12855_ ( .A(_09367_ ), .B(\pc_out[12] ), .Z(_09368_ ) );
AOI22_X1 _12856_ ( .A1(\alu_result_out[12] ), .A2(_09290_ ), .B1(_09291_ ), .B2(_09368_ ), .ZN(_09369_ ) );
NOR2_X1 _12857_ ( .A1(_09369_ ), .A2(\u_ifu.reset_sync ), .ZN(_00120_ ) );
NAND2_X1 _12858_ ( .A1(_09029_ ), .A2(_09033_ ), .ZN(_09370_ ) );
AOI21_X1 _12859_ ( .A(_09215_ ), .B1(_09370_ ), .B2(_09217_ ), .ZN(_09371_ ) );
OR2_X1 _12860_ ( .A1(_09371_ ), .A2(_09220_ ), .ZN(_09372_ ) );
XNOR2_X1 _12861_ ( .A(_09372_ ), .B(_09212_ ), .ZN(\alu_result_out[11] ) );
NAND2_X1 _12862_ ( .A1(\alu_result_out[11] ), .A2(_09107_ ), .ZN(_09373_ ) );
INV_X1 _12863_ ( .A(dnpc_$_MUX__Y_21_A_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_09374_ ) );
AND3_X1 _12864_ ( .A1(_09000_ ), .A2(_09374_ ), .A3(_09296_ ), .ZN(_09375_ ) );
XNOR2_X1 _12865_ ( .A(_09375_ ), .B(\pc_out[11] ), .ZN(_09376_ ) );
OR2_X1 _12866_ ( .A1(jump_en ), .A2(_09376_ ), .ZN(_09377_ ) );
AOI21_X1 _12867_ ( .A(\u_ifu.reset_sync ), .B1(_09373_ ), .B2(_09377_ ), .ZN(_00121_ ) );
XOR2_X1 _12868_ ( .A(_09273_ ), .B(_09280_ ), .Z(\alu_result_out[28] ) );
XNOR2_X1 _12869_ ( .A(_09312_ ), .B(dnpc_$_MUX__Y_3_A_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_09378_ ) );
AOI22_X1 _12870_ ( .A1(\alu_result_out[28] ), .A2(_09290_ ), .B1(_09291_ ), .B2(_09378_ ), .ZN(_09379_ ) );
NOR2_X1 _12871_ ( .A1(_09379_ ), .A2(\u_ifu.reset_sync ), .ZN(_00122_ ) );
NAND2_X1 _12872_ ( .A1(_09370_ ), .A2(_09217_ ), .ZN(_09380_ ) );
XNOR2_X1 _12873_ ( .A(_09380_ ), .B(_09215_ ), .ZN(\alu_result_out[10] ) );
NAND2_X1 _12874_ ( .A1(\alu_result_out[10] ), .A2(_09107_ ), .ZN(_09381_ ) );
AOI21_X1 _12875_ ( .A(_09374_ ), .B1(_09000_ ), .B2(_09296_ ), .ZN(_09382_ ) );
OR3_X1 _12876_ ( .A1(jump_en ), .A2(_09375_ ), .A3(_09382_ ), .ZN(_09383_ ) );
AOI21_X1 _12877_ ( .A(\u_ifu.reset_sync ), .B1(_09381_ ), .B2(_09383_ ), .ZN(_00123_ ) );
AOI21_X1 _12878_ ( .A(\u_ifu.reset_sync ), .B1(_09037_ ), .B2(_09041_ ), .ZN(_00124_ ) );
AND3_X1 _12879_ ( .A1(_09021_ ), .A2(_09098_ ), .A3(_09024_ ), .ZN(_00125_ ) );
AND3_X1 _12880_ ( .A1(_08998_ ), .A2(_09098_ ), .A3(_09004_ ), .ZN(_00126_ ) );
AOI21_X1 _12881_ ( .A(\u_ifu.reset_sync ), .B1(_09047_ ), .B2(_09049_ ), .ZN(_00127_ ) );
AND3_X1 _12882_ ( .A1(_09057_ ), .A2(_09098_ ), .A3(_09062_ ), .ZN(_00128_ ) );
AND2_X1 _12883_ ( .A1(_09075_ ), .A2(_09098_ ), .ZN(_00130_ ) );
INV_X1 _12884_ ( .A(_09256_ ), .ZN(_09384_ ) );
NAND2_X1 _12885_ ( .A1(_09250_ ), .A2(_09263_ ), .ZN(_09385_ ) );
AOI21_X1 _12886_ ( .A(_09384_ ), .B1(_09385_ ), .B2(_09269_ ), .ZN(_09386_ ) );
NOR2_X1 _12887_ ( .A1(_09386_ ), .A2(_09265_ ), .ZN(_09387_ ) );
XNOR2_X1 _12888_ ( .A(_09387_ ), .B(_09253_ ), .ZN(\alu_result_out[27] ) );
NAND2_X1 _12889_ ( .A1(\alu_result_out[27] ), .A2(_09107_ ), .ZN(_09388_ ) );
INV_X1 _12890_ ( .A(dnpc_$_MUX__Y_5_A_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_09389_ ) );
AND3_X1 _12891_ ( .A1(_09298_ ), .A2(_09389_ ), .A3(_09302_ ), .ZN(_09390_ ) );
XNOR2_X1 _12892_ ( .A(_09390_ ), .B(\pc_out[27] ), .ZN(_09391_ ) );
OR2_X1 _12893_ ( .A1(jump_en ), .A2(_09391_ ), .ZN(_09392_ ) );
AOI21_X1 _12894_ ( .A(\u_ifu.reset_sync ), .B1(_09388_ ), .B2(_09392_ ), .ZN(_00132_ ) );
AOI21_X1 _12895_ ( .A(_09270_ ), .B1(_09250_ ), .B2(_09263_ ), .ZN(_09393_ ) );
XNOR2_X1 _12896_ ( .A(_09393_ ), .B(_09256_ ), .ZN(\alu_result_out[26] ) );
XNOR2_X1 _12897_ ( .A(_09311_ ), .B(dnpc_$_MUX__Y_5_A_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_09394_ ) );
AOI22_X1 _12898_ ( .A1(\alu_result_out[26] ), .A2(_09290_ ), .B1(_09291_ ), .B2(_09394_ ), .ZN(_09395_ ) );
NOR2_X1 _12899_ ( .A1(_09395_ ), .A2(\u_ifu.reset_sync ), .ZN(_00133_ ) );
AND2_X1 _12900_ ( .A1(_09250_ ), .A2(_09259_ ), .ZN(_09396_ ) );
NOR2_X1 _12901_ ( .A1(_09396_ ), .A2(_09267_ ), .ZN(_09397_ ) );
XNOR2_X1 _12902_ ( .A(_09397_ ), .B(_09262_ ), .ZN(\alu_result_out[25] ) );
AND3_X1 _12903_ ( .A1(_09363_ ), .A2(\pc_out[13] ), .A3(_09294_ ), .ZN(_09398_ ) );
AND3_X1 _12904_ ( .A1(_09398_ ), .A2(\pc_out[17] ), .A3(\pc_out[16] ), .ZN(_09399_ ) );
AND2_X1 _12905_ ( .A1(_09399_ ), .A2(_09299_ ), .ZN(_09400_ ) );
AND3_X1 _12906_ ( .A1(_09400_ ), .A2(\pc_out[21] ), .A3(\pc_out[20] ), .ZN(_09401_ ) );
AND3_X1 _12907_ ( .A1(_09401_ ), .A2(\pc_out[24] ), .A3(_09301_ ), .ZN(_09402_ ) );
XOR2_X1 _12908_ ( .A(_09402_ ), .B(\pc_out[25] ), .Z(_09403_ ) );
AOI22_X1 _12909_ ( .A1(\alu_result_out[25] ), .A2(_09290_ ), .B1(_09291_ ), .B2(_09403_ ), .ZN(_09404_ ) );
NOR2_X1 _12910_ ( .A1(_09404_ ), .A2(\u_ifu.reset_sync ), .ZN(_00134_ ) );
XOR2_X1 _12911_ ( .A(_09250_ ), .B(_09259_ ), .Z(\alu_result_out[24] ) );
AND3_X1 _12912_ ( .A1(_09295_ ), .A2(_09297_ ), .A3(_09300_ ), .ZN(_09405_ ) );
AND2_X1 _12913_ ( .A1(_09405_ ), .A2(_09301_ ), .ZN(_09406_ ) );
XOR2_X1 _12914_ ( .A(_09406_ ), .B(\pc_out[24] ), .Z(_09407_ ) );
AOI22_X1 _12915_ ( .A1(\alu_result_out[24] ), .A2(_09036_ ), .B1(_08930_ ), .B2(_09407_ ), .ZN(_09408_ ) );
NOR2_X1 _12916_ ( .A1(_09408_ ), .A2(\u_ifu.reset_sync ), .ZN(_00135_ ) );
AOI21_X1 _12917_ ( .A(_09191_ ), .B1(_09317_ ), .B2(_09173_ ), .ZN(_09409_ ) );
AOI21_X1 _12918_ ( .A(_09196_ ), .B1(_09409_ ), .B2(_09186_ ), .ZN(_09410_ ) );
NOR2_X1 _12919_ ( .A1(_09410_ ), .A2(_09181_ ), .ZN(_09411_ ) );
NOR2_X1 _12920_ ( .A1(_09179_ ), .A2(_09180_ ), .ZN(_09412_ ) );
OR2_X1 _12921_ ( .A1(_09411_ ), .A2(_09412_ ), .ZN(_09413_ ) );
XNOR2_X1 _12922_ ( .A(_09413_ ), .B(_09177_ ), .ZN(\alu_result_out[23] ) );
NAND2_X1 _12923_ ( .A1(\alu_result_out[23] ), .A2(_09107_ ), .ZN(_09414_ ) );
INV_X1 _12924_ ( .A(_09405_ ), .ZN(_09415_ ) );
NOR2_X1 _12925_ ( .A1(_09415_ ), .A2(dnpc_$_MUX__Y_9_A_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_09416_ ) );
XNOR2_X1 _12926_ ( .A(_09416_ ), .B(\pc_out[23] ), .ZN(_09417_ ) );
OR2_X1 _12927_ ( .A1(jump_en ), .A2(_09417_ ), .ZN(_09418_ ) );
AOI21_X1 _12928_ ( .A(\u_ifu.reset_sync ), .B1(_09414_ ), .B2(_09418_ ), .ZN(_00136_ ) );
XOR2_X1 _12929_ ( .A(_09410_ ), .B(_09181_ ), .Z(\alu_result_out[22] ) );
XNOR2_X1 _12930_ ( .A(_09405_ ), .B(dnpc_$_MUX__Y_9_A_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_09419_ ) );
AOI22_X1 _12931_ ( .A1(\alu_result_out[22] ), .A2(_09036_ ), .B1(_08930_ ), .B2(_09419_ ), .ZN(_09420_ ) );
NOR2_X1 _12932_ ( .A1(_09420_ ), .A2(\u_ifu.reset_sync ), .ZN(_00137_ ) );
INV_X1 _12933_ ( .A(_09409_ ), .ZN(_09421_ ) );
NAND2_X1 _12934_ ( .A1(_09421_ ), .A2(_09195_ ), .ZN(_09422_ ) );
XNOR2_X1 _12935_ ( .A(_09422_ ), .B(_09187_ ), .ZN(\alu_result_out[21] ) );
NAND2_X1 _12936_ ( .A1(\alu_result_out[21] ), .A2(_09107_ ), .ZN(_09423_ ) );
NOR2_X1 _12937_ ( .A1(_09319_ ), .A2(dnpc_$_MUX__Y_11_A_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_09424_ ) );
XNOR2_X1 _12938_ ( .A(_09424_ ), .B(\pc_out[21] ), .ZN(_09425_ ) );
OR2_X1 _12939_ ( .A1(jump_en ), .A2(_09425_ ), .ZN(_09426_ ) );
AOI21_X1 _12940_ ( .A(\u_ifu.reset_sync ), .B1(_09423_ ), .B2(_09426_ ), .ZN(_00138_ ) );
INV_X1 _12941_ ( .A(_09304_ ), .ZN(_09427_ ) );
OR2_X1 _12942_ ( .A1(_09427_ ), .A2(dnpc_$_MUX__Y_1_A_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_09428_ ) );
XNOR2_X1 _12943_ ( .A(_09428_ ), .B(\pc_out[31] ), .ZN(_09429_ ) );
NAND3_X1 _12944_ ( .A1(_08906_ ), .A2(_08929_ ), .A3(_09429_ ), .ZN(_09430_ ) );
OR2_X1 _12945_ ( .A1(_09284_ ), .A2(_09289_ ), .ZN(_09431_ ) );
NAND3_X1 _12946_ ( .A1(_09288_ ), .A2(_08856_ ), .A3(_09175_ ), .ZN(_09432_ ) );
NAND2_X1 _12947_ ( .A1(_09431_ ), .A2(_09432_ ), .ZN(_09433_ ) );
NOR2_X1 _12948_ ( .A1(_08953_ ), .A2(_08837_ ), .ZN(_09434_ ) );
NAND3_X1 _12949_ ( .A1(_08832_ ), .A2(_08611_ ), .A3(_08997_ ), .ZN(_09435_ ) );
NAND3_X1 _12950_ ( .A1(_08905_ ), .A2(\ifu_rdata[0] ), .A3(\pc_out[31] ), .ZN(_09436_ ) );
AND2_X1 _12951_ ( .A1(_09435_ ), .A2(_09436_ ), .ZN(_09437_ ) );
XNOR2_X1 _12952_ ( .A(_09434_ ), .B(_09437_ ), .ZN(_09438_ ) );
XOR2_X1 _12953_ ( .A(_09433_ ), .B(_09438_ ), .Z(\alu_result_out[31] ) );
INV_X1 _12954_ ( .A(\alu_result_out[31] ), .ZN(_09439_ ) );
OAI211_X1 _12955_ ( .A(_09098_ ), .B(_09430_ ), .C1(_09439_ ), .C2(_09087_ ), .ZN(_00139_ ) );
INV_X1 _12956_ ( .A(_09136_ ), .ZN(_09440_ ) );
BUF_X4 _12957_ ( .A(_09440_ ), .Z(_09441_ ) );
INV_X8 _12958_ ( .A(_09140_ ), .ZN(_09442_ ) );
BUF_X8 _12959_ ( .A(_09442_ ), .Z(_09443_ ) );
BUF_X4 _12960_ ( .A(_09443_ ), .Z(_09444_ ) );
OAI21_X1 _12961_ ( .A(\u_lsu.pmem[4387] ), .B1(_09441_ ), .B2(_09444_ ), .ZN(_09445_ ) );
INV_X1 _12962_ ( .A(_08650_ ), .ZN(_09446_ ) );
NOR2_X4 _12963_ ( .A1(_09145_ ), .A2(_09446_ ), .ZN(_09447_ ) );
BUF_X4 _12964_ ( .A(_09447_ ), .Z(_09448_ ) );
BUF_X4 _12965_ ( .A(_09448_ ), .Z(_09449_ ) );
BUF_X8 _12966_ ( .A(_09140_ ), .Z(_09450_ ) );
BUF_X8 _12967_ ( .A(_09450_ ), .Z(_09451_ ) );
BUF_X4 _12968_ ( .A(_09451_ ), .Z(_09452_ ) );
INV_X4 _12969_ ( .A(_09134_ ), .ZN(_09453_ ) );
BUF_X4 _12970_ ( .A(_09453_ ), .Z(_09454_ ) );
BUF_X8 _12971_ ( .A(_09454_ ), .Z(_09455_ ) );
BUF_X4 _12972_ ( .A(_09455_ ), .Z(_09456_ ) );
NAND4_X1 _12973_ ( .A1(_09449_ ), .A2(_09452_ ), .A3(_09131_ ), .A4(_09456_ ), .ZN(_09457_ ) );
AOI21_X1 _12974_ ( .A(fanout_net_8 ), .B1(_09445_ ), .B2(_09457_ ), .ZN(_00140_ ) );
BUF_X16 _12975_ ( .A(_09442_ ), .Z(_09458_ ) );
BUF_X8 _12976_ ( .A(_09458_ ), .Z(_09459_ ) );
BUF_X4 _12977_ ( .A(_09459_ ), .Z(_09460_ ) );
BUF_X4 _12978_ ( .A(_09453_ ), .Z(_09461_ ) );
BUF_X4 _12979_ ( .A(_09130_ ), .Z(_09462_ ) );
BUF_X2 _12980_ ( .A(_09054_ ), .Z(_09463_ ) );
INV_X1 _12981_ ( .A(_09113_ ), .ZN(_09464_ ) );
NOR2_X1 _12982_ ( .A1(_09463_ ), .A2(_09464_ ), .ZN(_09465_ ) );
INV_X1 _12983_ ( .A(_09465_ ), .ZN(_09466_ ) );
NOR3_X2 _12984_ ( .A1(_09118_ ), .A2(_09462_ ), .A3(_09466_ ), .ZN(_09467_ ) );
NAND2_X1 _12985_ ( .A1(_09461_ ), .A2(_09467_ ), .ZN(_09468_ ) );
BUF_X4 _12986_ ( .A(_09468_ ), .Z(_09469_ ) );
OAI21_X1 _12987_ ( .A(\u_lsu.pmem[4354] ), .B1(_09460_ ), .B2(_09469_ ), .ZN(_09470_ ) );
BUF_X16 _12988_ ( .A(_09140_ ), .Z(_09471_ ) );
BUF_X8 _12989_ ( .A(_09471_ ), .Z(_09472_ ) );
BUF_X4 _12990_ ( .A(_09472_ ), .Z(_09473_ ) );
BUF_X4 _12991_ ( .A(_08659_ ), .Z(_09474_ ) );
BUF_X4 _12992_ ( .A(_09453_ ), .Z(_09475_ ) );
BUF_X8 _12993_ ( .A(_09475_ ), .Z(_09476_ ) );
BUF_X4 _12994_ ( .A(_09476_ ), .Z(_09477_ ) );
NAND4_X1 _12995_ ( .A1(_09473_ ), .A2(_09474_ ), .A3(_09477_ ), .A4(_09467_ ), .ZN(_09478_ ) );
AOI21_X1 _12996_ ( .A(fanout_net_8 ), .B1(_09470_ ), .B2(_09478_ ), .ZN(_00141_ ) );
INV_X1 _12997_ ( .A(_09053_ ), .ZN(_09479_ ) );
BUF_X4 _12998_ ( .A(_09479_ ), .Z(_09480_ ) );
BUF_X8 _12999_ ( .A(_09480_ ), .Z(_09481_ ) );
BUF_X4 _13000_ ( .A(_09481_ ), .Z(_09482_ ) );
BUF_X4 _13001_ ( .A(_09083_ ), .Z(_09483_ ) );
BUF_X4 _13002_ ( .A(_09123_ ), .Z(_09484_ ) );
AND2_X2 _13003_ ( .A1(_09483_ ), .A2(_09484_ ), .ZN(_09485_ ) );
AND2_X1 _13004_ ( .A1(_09482_ ), .A2(_09485_ ), .ZN(_09486_ ) );
BUF_X2 _13005_ ( .A(_09046_ ), .Z(_09487_ ) );
AND2_X1 _13006_ ( .A1(_09486_ ), .A2(_09487_ ), .ZN(_09488_ ) );
BUF_X2 _13007_ ( .A(_08993_ ), .Z(_09489_ ) );
AND2_X1 _13008_ ( .A1(_09488_ ), .A2(_09489_ ), .ZN(_09490_ ) );
CLKBUF_X2 _13009_ ( .A(_09018_ ), .Z(_09491_ ) );
AND2_X1 _13010_ ( .A1(_09490_ ), .A2(_09491_ ), .ZN(_09492_ ) );
BUF_X4 _13011_ ( .A(_09138_ ), .Z(_09493_ ) );
AND2_X1 _13012_ ( .A1(_09492_ ), .A2(_09493_ ), .ZN(_09494_ ) );
OAI21_X1 _13013_ ( .A(_09110_ ), .B1(_09494_ ), .B2(\u_lsu.pmem[4000] ), .ZN(_09495_ ) );
BUF_X4 _13014_ ( .A(_09493_ ), .Z(_09496_ ) );
CLKBUF_X2 _13015_ ( .A(_08952_ ), .Z(_09497_ ) );
CLKBUF_X2 _13016_ ( .A(_09137_ ), .Z(_09498_ ) );
CLKBUF_X2 _13017_ ( .A(_09498_ ), .Z(_09499_ ) );
OAI211_X1 _13018_ ( .A(_09492_ ), .B(_09496_ ), .C1(_09497_ ), .C2(_09499_ ), .ZN(_09500_ ) );
INV_X1 _13019_ ( .A(_09500_ ), .ZN(_09501_ ) );
NOR2_X1 _13020_ ( .A1(_09495_ ), .A2(_09501_ ), .ZN(_00142_ ) );
NOR2_X4 _13021_ ( .A1(_09144_ ), .A2(_09112_ ), .ZN(_09502_ ) );
AND2_X4 _13022_ ( .A1(_09502_ ), .A2(_09483_ ), .ZN(_09503_ ) );
AND2_X4 _13023_ ( .A1(_09503_ ), .A2(_09482_ ), .ZN(_09504_ ) );
BUF_X2 _13024_ ( .A(_09129_ ), .Z(_09505_ ) );
INV_X2 _13025_ ( .A(_09117_ ), .ZN(_09506_ ) );
AND3_X1 _13026_ ( .A1(_09504_ ), .A2(_09505_ ), .A3(_09506_ ), .ZN(_09507_ ) );
NAND2_X1 _13027_ ( .A1(_09507_ ), .A2(_09475_ ), .ZN(_09508_ ) );
BUF_X4 _13028_ ( .A(_09508_ ), .Z(_09509_ ) );
BUF_X4 _13029_ ( .A(_09472_ ), .Z(_09510_ ) );
OAI21_X1 _13030_ ( .A(\u_lsu.pmem[388] ), .B1(_09509_ ), .B2(_09510_ ), .ZN(_09511_ ) );
BUF_X4 _13031_ ( .A(_09507_ ), .Z(_09512_ ) );
BUF_X4 _13032_ ( .A(_09512_ ), .Z(_09513_ ) );
BUF_X4 _13033_ ( .A(_08605_ ), .Z(_09514_ ) );
BUF_X8 _13034_ ( .A(_09442_ ), .Z(_09515_ ) );
BUF_X4 _13035_ ( .A(_09515_ ), .Z(_09516_ ) );
NAND4_X1 _13036_ ( .A1(_09513_ ), .A2(_09514_ ), .A3(_09477_ ), .A4(_09516_ ), .ZN(_09517_ ) );
AOI21_X1 _13037_ ( .A(fanout_net_8 ), .B1(_09511_ ), .B2(_09517_ ), .ZN(_00143_ ) );
OAI21_X1 _13038_ ( .A(\u_lsu.pmem[387] ), .B1(_09509_ ), .B2(_09510_ ), .ZN(_09518_ ) );
BUF_X4 _13039_ ( .A(_08650_ ), .Z(_09519_ ) );
BUF_X4 _13040_ ( .A(_09519_ ), .Z(_09520_ ) );
BUF_X4 _13041_ ( .A(_09476_ ), .Z(_09521_ ) );
BUF_X8 _13042_ ( .A(_09442_ ), .Z(_09522_ ) );
BUF_X4 _13043_ ( .A(_09522_ ), .Z(_09523_ ) );
NAND4_X1 _13044_ ( .A1(_09513_ ), .A2(_09520_ ), .A3(_09521_ ), .A4(_09523_ ), .ZN(_09524_ ) );
AOI21_X1 _13045_ ( .A(fanout_net_8 ), .B1(_09518_ ), .B2(_09524_ ), .ZN(_00144_ ) );
OAI21_X1 _13046_ ( .A(\u_lsu.pmem[386] ), .B1(_09509_ ), .B2(_09510_ ), .ZN(_09525_ ) );
BUF_X4 _13047_ ( .A(_09111_ ), .Z(_09526_ ) );
BUF_X4 _13048_ ( .A(_09526_ ), .Z(_09527_ ) );
BUF_X4 _13049_ ( .A(_09527_ ), .Z(_09528_ ) );
BUF_X4 _13050_ ( .A(_09528_ ), .Z(_09529_ ) );
BUF_X4 _13051_ ( .A(_09529_ ), .Z(_09530_ ) );
BUF_X4 _13052_ ( .A(_09530_ ), .Z(_09531_ ) );
XNOR2_X1 _13053_ ( .A(\alu_result_out[4] ), .B(_09531_ ), .ZN(_09532_ ) );
NAND3_X1 _13054_ ( .A1(_09502_ ), .A2(_08659_ ), .A3(_09532_ ), .ZN(_09533_ ) );
XNOR2_X1 _13055_ ( .A(_09054_ ), .B(_09464_ ), .ZN(_09534_ ) );
BUF_X2 _13056_ ( .A(_09534_ ), .Z(_09535_ ) );
BUF_X4 _13057_ ( .A(_09462_ ), .Z(_09536_ ) );
NOR3_X1 _13058_ ( .A1(_09533_ ), .A2(_09535_ ), .A3(_09536_ ), .ZN(_09537_ ) );
BUF_X4 _13059_ ( .A(_09506_ ), .Z(_09538_ ) );
BUF_X8 _13060_ ( .A(_09538_ ), .Z(_09539_ ) );
BUF_X4 _13061_ ( .A(_09539_ ), .Z(_09540_ ) );
NAND4_X1 _13062_ ( .A1(_09537_ ), .A2(_09540_ ), .A3(_09521_ ), .A4(_09523_ ), .ZN(_09541_ ) );
AOI21_X1 _13063_ ( .A(fanout_net_8 ), .B1(_09525_ ), .B2(_09541_ ), .ZN(_00145_ ) );
OAI21_X1 _13064_ ( .A(\u_lsu.pmem[385] ), .B1(_09509_ ), .B2(_09510_ ), .ZN(_09542_ ) );
BUF_X4 _13065_ ( .A(_08638_ ), .Z(_09543_ ) );
BUF_X4 _13066_ ( .A(_09543_ ), .Z(_09544_ ) );
NAND4_X1 _13067_ ( .A1(_09513_ ), .A2(_09544_ ), .A3(_09521_ ), .A4(_09523_ ), .ZN(_09545_ ) );
AOI21_X1 _13068_ ( .A(fanout_net_8 ), .B1(_09542_ ), .B2(_09545_ ), .ZN(_00146_ ) );
OAI21_X1 _13069_ ( .A(\u_lsu.pmem[384] ), .B1(_09509_ ), .B2(_09510_ ), .ZN(_09546_ ) );
BUF_X4 _13070_ ( .A(_08631_ ), .Z(_09547_ ) );
BUF_X4 _13071_ ( .A(_09547_ ), .Z(_09548_ ) );
NAND4_X1 _13072_ ( .A1(_09513_ ), .A2(_09548_ ), .A3(_09521_ ), .A4(_09523_ ), .ZN(_09549_ ) );
AOI21_X1 _13073_ ( .A(fanout_net_8 ), .B1(_09546_ ), .B2(_09549_ ), .ZN(_00147_ ) );
BUF_X4 _13074_ ( .A(_09054_ ), .Z(_09550_ ) );
AND2_X4 _13075_ ( .A1(_09066_ ), .A2(_09089_ ), .ZN(_09551_ ) );
BUF_X16 _13076_ ( .A(_09551_ ), .Z(_09552_ ) );
BUF_X16 _13077_ ( .A(_09552_ ), .Z(_09553_ ) );
BUF_X32 _13078_ ( .A(_09553_ ), .Z(_09554_ ) );
INV_X1 _13079_ ( .A(_09554_ ), .ZN(_09555_ ) );
NOR2_X4 _13080_ ( .A1(_09555_ ), .A2(_09083_ ), .ZN(_09556_ ) );
INV_X1 _13081_ ( .A(_09556_ ), .ZN(_09557_ ) );
NOR3_X2 _13082_ ( .A1(_09046_ ), .A2(_09550_ ), .A3(_09557_ ), .ZN(_09558_ ) );
INV_X1 _13083_ ( .A(_09558_ ), .ZN(_09559_ ) );
NOR3_X4 _13084_ ( .A1(_09134_ ), .A2(_09118_ ), .A3(_09559_ ), .ZN(_09560_ ) );
INV_X1 _13085_ ( .A(_09560_ ), .ZN(_09561_ ) );
BUF_X8 _13086_ ( .A(_09141_ ), .Z(_09562_ ) );
NOR2_X2 _13087_ ( .A1(_09561_ ), .A2(_09562_ ), .ZN(_09563_ ) );
OAI21_X1 _13088_ ( .A(_09110_ ), .B1(_09563_ ), .B2(\u_lsu.pmem[359] ), .ZN(_09564_ ) );
INV_X1 _13089_ ( .A(_08582_ ), .ZN(_09565_ ) );
NOR2_X4 _13090_ ( .A1(_09144_ ), .A2(_09565_ ), .ZN(_09566_ ) );
INV_X1 _13091_ ( .A(_09566_ ), .ZN(_09567_ ) );
BUF_X4 _13092_ ( .A(_09567_ ), .Z(_09568_ ) );
AOI21_X1 _13093_ ( .A(_09564_ ), .B1(_09563_ ), .B2(_09568_ ), .ZN(_00148_ ) );
BUF_X4 _13094_ ( .A(_09561_ ), .Z(_09569_ ) );
BUF_X4 _13095_ ( .A(_09472_ ), .Z(_09570_ ) );
OAI21_X1 _13096_ ( .A(\u_lsu.pmem[358] ), .B1(_09569_ ), .B2(_09570_ ), .ZN(_09571_ ) );
BUF_X8 _13097_ ( .A(_09458_ ), .Z(_09572_ ) );
BUF_X4 _13098_ ( .A(_09572_ ), .Z(_09573_ ) );
BUF_X4 _13099_ ( .A(_09560_ ), .Z(_09574_ ) );
BUF_X4 _13100_ ( .A(_08617_ ), .Z(_09575_ ) );
INV_X1 _13101_ ( .A(_09575_ ), .ZN(_09576_ ) );
NOR2_X4 _13102_ ( .A1(_09144_ ), .A2(_09576_ ), .ZN(_09577_ ) );
BUF_X4 _13103_ ( .A(_09577_ ), .Z(_09578_ ) );
BUF_X4 _13104_ ( .A(_09578_ ), .Z(_09579_ ) );
NAND3_X1 _13105_ ( .A1(_09573_ ), .A2(_09574_ ), .A3(_09579_ ), .ZN(_09580_ ) );
AOI21_X1 _13106_ ( .A(fanout_net_8 ), .B1(_09571_ ), .B2(_09580_ ), .ZN(_00149_ ) );
OAI21_X1 _13107_ ( .A(\u_lsu.pmem[357] ), .B1(_09569_ ), .B2(_09570_ ), .ZN(_09581_ ) );
BUF_X4 _13108_ ( .A(_08595_ ), .Z(_09582_ ) );
INV_X1 _13109_ ( .A(_09582_ ), .ZN(_09583_ ) );
NOR2_X4 _13110_ ( .A1(_09144_ ), .A2(_09583_ ), .ZN(_09584_ ) );
BUF_X4 _13111_ ( .A(_09584_ ), .Z(_09585_ ) );
BUF_X4 _13112_ ( .A(_09585_ ), .Z(_09586_ ) );
NAND3_X1 _13113_ ( .A1(_09573_ ), .A2(_09574_ ), .A3(_09586_ ), .ZN(_09587_ ) );
AOI21_X1 _13114_ ( .A(fanout_net_8 ), .B1(_09581_ ), .B2(_09587_ ), .ZN(_00150_ ) );
OAI21_X1 _13115_ ( .A(\u_lsu.pmem[356] ), .B1(_09569_ ), .B2(_09570_ ), .ZN(_09588_ ) );
BUF_X4 _13116_ ( .A(_09148_ ), .Z(_09589_ ) );
NAND3_X1 _13117_ ( .A1(_09573_ ), .A2(_09589_ ), .A3(_09560_ ), .ZN(_09590_ ) );
AOI21_X1 _13118_ ( .A(fanout_net_8 ), .B1(_09588_ ), .B2(_09590_ ), .ZN(_00151_ ) );
OAI21_X1 _13119_ ( .A(\u_lsu.pmem[355] ), .B1(_09569_ ), .B2(_09570_ ), .ZN(_09591_ ) );
BUF_X4 _13120_ ( .A(_09448_ ), .Z(_09592_ ) );
NAND3_X1 _13121_ ( .A1(_09573_ ), .A2(_09592_ ), .A3(_09560_ ), .ZN(_09593_ ) );
AOI21_X1 _13122_ ( .A(fanout_net_8 ), .B1(_09591_ ), .B2(_09593_ ), .ZN(_00152_ ) );
BUF_X2 _13123_ ( .A(_09046_ ), .Z(_09594_ ) );
AND2_X4 _13124_ ( .A1(_09504_ ), .A2(_09594_ ), .ZN(_09595_ ) );
AND2_X4 _13125_ ( .A1(_09595_ ), .A2(_09489_ ), .ZN(_09596_ ) );
AND2_X4 _13126_ ( .A1(_09596_ ), .A2(_09491_ ), .ZN(_09597_ ) );
INV_X8 _13127_ ( .A(_09597_ ), .ZN(_09598_ ) );
BUF_X8 _13128_ ( .A(_09598_ ), .Z(_09599_ ) );
OAI21_X1 _13129_ ( .A(\u_lsu.pmem[3975] ), .B1(_09599_ ), .B2(_09570_ ), .ZN(_09600_ ) );
BUF_X4 _13130_ ( .A(_09596_ ), .Z(_09601_ ) );
BUF_X4 _13131_ ( .A(_09601_ ), .Z(_09602_ ) );
BUF_X4 _13132_ ( .A(_08582_ ), .Z(_09603_ ) );
BUF_X4 _13133_ ( .A(_09018_ ), .Z(_09604_ ) );
BUF_X4 _13134_ ( .A(_09604_ ), .Z(_09605_ ) );
BUF_X4 _13135_ ( .A(_09605_ ), .Z(_09606_ ) );
BUF_X4 _13136_ ( .A(_09606_ ), .Z(_09607_ ) );
NAND4_X1 _13137_ ( .A1(_09602_ ), .A2(_09603_ ), .A3(_09607_ ), .A4(_09523_ ), .ZN(_09608_ ) );
AOI21_X1 _13138_ ( .A(fanout_net_8 ), .B1(_09600_ ), .B2(_09608_ ), .ZN(_00153_ ) );
OAI21_X1 _13139_ ( .A(\u_lsu.pmem[354] ), .B1(_09569_ ), .B2(_09570_ ), .ZN(_09609_ ) );
NOR2_X4 _13140_ ( .A1(_09145_ ), .A2(_08962_ ), .ZN(_09610_ ) );
BUF_X4 _13141_ ( .A(_09610_ ), .Z(_09611_ ) );
BUF_X4 _13142_ ( .A(_09611_ ), .Z(_09612_ ) );
NAND3_X1 _13143_ ( .A1(_09573_ ), .A2(_09612_ ), .A3(_09560_ ), .ZN(_09613_ ) );
AOI21_X1 _13144_ ( .A(fanout_net_8 ), .B1(_09609_ ), .B2(_09613_ ), .ZN(_00154_ ) );
OAI21_X1 _13145_ ( .A(\u_lsu.pmem[353] ), .B1(_09569_ ), .B2(_09570_ ), .ZN(_09614_ ) );
NOR2_X1 _13146_ ( .A1(_09145_ ), .A2(_08639_ ), .ZN(_09615_ ) );
BUF_X4 _13147_ ( .A(_09615_ ), .Z(_09616_ ) );
BUF_X4 _13148_ ( .A(_09616_ ), .Z(_09617_ ) );
NAND3_X1 _13149_ ( .A1(_09573_ ), .A2(_09617_ ), .A3(_09560_ ), .ZN(_09618_ ) );
AOI21_X1 _13150_ ( .A(fanout_net_8 ), .B1(_09614_ ), .B2(_09618_ ), .ZN(_00155_ ) );
OAI21_X1 _13151_ ( .A(\u_lsu.pmem[352] ), .B1(_09569_ ), .B2(_09570_ ), .ZN(_09619_ ) );
NOR2_X4 _13152_ ( .A1(_09144_ ), .A2(_08952_ ), .ZN(_09620_ ) );
BUF_X4 _13153_ ( .A(_09620_ ), .Z(_09621_ ) );
BUF_X4 _13154_ ( .A(_09621_ ), .Z(_09622_ ) );
NAND3_X1 _13155_ ( .A1(_09573_ ), .A2(_09622_ ), .A3(_09560_ ), .ZN(_09623_ ) );
AOI21_X1 _13156_ ( .A(fanout_net_8 ), .B1(_09619_ ), .B2(_09623_ ), .ZN(_00156_ ) );
AND2_X4 _13157_ ( .A1(_09066_ ), .A2(_09090_ ), .ZN(_09624_ ) );
BUF_X4 _13158_ ( .A(_09624_ ), .Z(_09625_ ) );
BUF_X16 _13159_ ( .A(_09625_ ), .Z(_09626_ ) );
BUF_X16 _13160_ ( .A(_09626_ ), .Z(_09627_ ) );
INV_X1 _13161_ ( .A(_09627_ ), .ZN(_09628_ ) );
NOR2_X2 _13162_ ( .A1(_09628_ ), .A2(_09083_ ), .ZN(_09629_ ) );
INV_X1 _13163_ ( .A(_09629_ ), .ZN(_09630_ ) );
NOR3_X1 _13164_ ( .A1(_09046_ ), .A2(_09550_ ), .A3(_09630_ ), .ZN(_09631_ ) );
INV_X1 _13165_ ( .A(_09631_ ), .ZN(_09632_ ) );
NOR3_X4 _13166_ ( .A1(_09134_ ), .A2(_09118_ ), .A3(_09632_ ), .ZN(_09633_ ) );
INV_X1 _13167_ ( .A(_09633_ ), .ZN(_09634_ ) );
BUF_X4 _13168_ ( .A(_09471_ ), .Z(_09635_ ) );
NOR2_X1 _13169_ ( .A1(_09634_ ), .A2(_09635_ ), .ZN(_09636_ ) );
OAI21_X1 _13170_ ( .A(_09110_ ), .B1(_09636_ ), .B2(\u_lsu.pmem[327] ), .ZN(_09637_ ) );
BUF_X4 _13171_ ( .A(_09567_ ), .Z(_09638_ ) );
AOI21_X1 _13172_ ( .A(_09637_ ), .B1(_09638_ ), .B2(_09636_ ), .ZN(_00157_ ) );
BUF_X4 _13173_ ( .A(_09634_ ), .Z(_09639_ ) );
OAI21_X1 _13174_ ( .A(\u_lsu.pmem[326] ), .B1(_09639_ ), .B2(_09570_ ), .ZN(_09640_ ) );
BUF_X8 _13175_ ( .A(_09458_ ), .Z(_09641_ ) );
BUF_X4 _13176_ ( .A(_09641_ ), .Z(_09642_ ) );
BUF_X4 _13177_ ( .A(_09633_ ), .Z(_09643_ ) );
NAND3_X1 _13178_ ( .A1(_09642_ ), .A2(_09579_ ), .A3(_09643_ ), .ZN(_09644_ ) );
AOI21_X1 _13179_ ( .A(fanout_net_8 ), .B1(_09640_ ), .B2(_09644_ ), .ZN(_00158_ ) );
OAI21_X1 _13180_ ( .A(\u_lsu.pmem[325] ), .B1(_09639_ ), .B2(_09570_ ), .ZN(_09645_ ) );
NAND3_X1 _13181_ ( .A1(_09642_ ), .A2(_09586_ ), .A3(_09643_ ), .ZN(_09646_ ) );
AOI21_X1 _13182_ ( .A(fanout_net_8 ), .B1(_09645_ ), .B2(_09646_ ), .ZN(_00159_ ) );
BUF_X8 _13183_ ( .A(_09471_ ), .Z(_09647_ ) );
BUF_X4 _13184_ ( .A(_09647_ ), .Z(_09648_ ) );
OAI21_X1 _13185_ ( .A(\u_lsu.pmem[324] ), .B1(_09639_ ), .B2(_09648_ ), .ZN(_09649_ ) );
NAND3_X1 _13186_ ( .A1(_09642_ ), .A2(_09589_ ), .A3(_09633_ ), .ZN(_09650_ ) );
AOI21_X1 _13187_ ( .A(fanout_net_8 ), .B1(_09649_ ), .B2(_09650_ ), .ZN(_00160_ ) );
OAI21_X1 _13188_ ( .A(\u_lsu.pmem[323] ), .B1(_09639_ ), .B2(_09648_ ), .ZN(_09651_ ) );
NAND3_X1 _13189_ ( .A1(_09642_ ), .A2(_09592_ ), .A3(_09633_ ), .ZN(_09652_ ) );
AOI21_X1 _13190_ ( .A(fanout_net_8 ), .B1(_09651_ ), .B2(_09652_ ), .ZN(_00161_ ) );
OAI21_X1 _13191_ ( .A(\u_lsu.pmem[322] ), .B1(_09639_ ), .B2(_09648_ ), .ZN(_09653_ ) );
NAND3_X1 _13192_ ( .A1(_09642_ ), .A2(_09612_ ), .A3(_09633_ ), .ZN(_09654_ ) );
AOI21_X1 _13193_ ( .A(fanout_net_8 ), .B1(_09653_ ), .B2(_09654_ ), .ZN(_00162_ ) );
OAI21_X1 _13194_ ( .A(\u_lsu.pmem[321] ), .B1(_09639_ ), .B2(_09648_ ), .ZN(_09655_ ) );
NAND3_X1 _13195_ ( .A1(_09642_ ), .A2(_09617_ ), .A3(_09633_ ), .ZN(_09656_ ) );
AOI21_X1 _13196_ ( .A(fanout_net_8 ), .B1(_09655_ ), .B2(_09656_ ), .ZN(_00163_ ) );
OAI21_X1 _13197_ ( .A(\u_lsu.pmem[3974] ), .B1(_09599_ ), .B2(_09648_ ), .ZN(_09657_ ) );
BUF_X4 _13198_ ( .A(_09575_ ), .Z(_09658_ ) );
BUF_X4 _13199_ ( .A(_09606_ ), .Z(_09659_ ) );
NAND4_X1 _13200_ ( .A1(_09602_ ), .A2(_09658_ ), .A3(_09659_ ), .A4(_09523_ ), .ZN(_09660_ ) );
AOI21_X1 _13201_ ( .A(fanout_net_8 ), .B1(_09657_ ), .B2(_09660_ ), .ZN(_00164_ ) );
OAI21_X1 _13202_ ( .A(\u_lsu.pmem[320] ), .B1(_09639_ ), .B2(_09648_ ), .ZN(_09661_ ) );
NAND3_X1 _13203_ ( .A1(_09642_ ), .A2(_09622_ ), .A3(_09633_ ), .ZN(_09662_ ) );
AOI21_X1 _13204_ ( .A(fanout_net_8 ), .B1(_09661_ ), .B2(_09662_ ), .ZN(_00165_ ) );
AND2_X1 _13205_ ( .A1(_09566_ ), .A2(_09125_ ), .ZN(_09663_ ) );
BUF_X4 _13206_ ( .A(_09115_ ), .Z(_09664_ ) );
BUF_X4 _13207_ ( .A(_09664_ ), .Z(_09665_ ) );
BUF_X4 _13208_ ( .A(_09665_ ), .Z(_09666_ ) );
BUF_X4 _13209_ ( .A(_09666_ ), .Z(_09667_ ) );
INV_X1 _13210_ ( .A(_09534_ ), .ZN(_09668_ ) );
BUF_X4 _13211_ ( .A(_09668_ ), .Z(_09669_ ) );
AND3_X2 _13212_ ( .A1(_09663_ ), .A2(_09667_ ), .A3(_09669_ ), .ZN(_09670_ ) );
BUF_X8 _13213_ ( .A(_09539_ ), .Z(_09671_ ) );
BUF_X4 _13214_ ( .A(_09671_ ), .Z(_09672_ ) );
BUF_X8 _13215_ ( .A(_09455_ ), .Z(_09673_ ) );
BUF_X4 _13216_ ( .A(_09673_ ), .Z(_09674_ ) );
BUF_X8 _13217_ ( .A(_09442_ ), .Z(_09675_ ) );
BUF_X4 _13218_ ( .A(_09675_ ), .Z(_09676_ ) );
NAND4_X1 _13219_ ( .A1(_09670_ ), .A2(_09672_ ), .A3(_09674_ ), .A4(_09676_ ), .ZN(_09677_ ) );
BUF_X4 _13220_ ( .A(_09451_ ), .Z(_09678_ ) );
OAI21_X1 _13221_ ( .A(\u_lsu.pmem[295] ), .B1(_09441_ ), .B2(_09678_ ), .ZN(_09679_ ) );
AOI21_X1 _13222_ ( .A(fanout_net_8 ), .B1(_09677_ ), .B2(_09679_ ), .ZN(_00166_ ) );
AND2_X1 _13223_ ( .A1(_09577_ ), .A2(_09125_ ), .ZN(_09680_ ) );
AND3_X2 _13224_ ( .A1(_09680_ ), .A2(_09667_ ), .A3(_09669_ ), .ZN(_09681_ ) );
NAND4_X1 _13225_ ( .A1(_09681_ ), .A2(_09672_ ), .A3(_09674_ ), .A4(_09676_ ), .ZN(_09682_ ) );
OAI21_X1 _13226_ ( .A(\u_lsu.pmem[294] ), .B1(_09441_ ), .B2(_09678_ ), .ZN(_09683_ ) );
AOI21_X1 _13227_ ( .A(fanout_net_8 ), .B1(_09682_ ), .B2(_09683_ ), .ZN(_00167_ ) );
AND2_X1 _13228_ ( .A1(_09584_ ), .A2(_09125_ ), .ZN(_09684_ ) );
AND3_X2 _13229_ ( .A1(_09684_ ), .A2(_09667_ ), .A3(_09669_ ), .ZN(_09685_ ) );
BUF_X4 _13230_ ( .A(_09673_ ), .Z(_09686_ ) );
NAND4_X1 _13231_ ( .A1(_09685_ ), .A2(_09672_ ), .A3(_09686_ ), .A4(_09676_ ), .ZN(_09687_ ) );
OAI21_X1 _13232_ ( .A(\u_lsu.pmem[293] ), .B1(_09441_ ), .B2(_09678_ ), .ZN(_09688_ ) );
AOI21_X1 _13233_ ( .A(fanout_net_8 ), .B1(_09687_ ), .B2(_09688_ ), .ZN(_00168_ ) );
AND2_X1 _13234_ ( .A1(_09522_ ), .A2(_09136_ ), .ZN(_09689_ ) );
OAI21_X1 _13235_ ( .A(_09110_ ), .B1(_09689_ ), .B2(\u_lsu.pmem[292] ), .ZN(_09690_ ) );
BUF_X4 _13236_ ( .A(_09149_ ), .Z(_09691_ ) );
AOI21_X1 _13237_ ( .A(_09690_ ), .B1(_09691_ ), .B2(_09689_ ), .ZN(_00169_ ) );
OAI21_X1 _13238_ ( .A(\u_lsu.pmem[291] ), .B1(_09441_ ), .B2(_09648_ ), .ZN(_09692_ ) );
NAND3_X1 _13239_ ( .A1(_09642_ ), .A2(_09136_ ), .A3(_09449_ ), .ZN(_09693_ ) );
AOI21_X1 _13240_ ( .A(fanout_net_8 ), .B1(_09692_ ), .B2(_09693_ ), .ZN(_00170_ ) );
OAI21_X1 _13241_ ( .A(\u_lsu.pmem[290] ), .B1(_09441_ ), .B2(_09648_ ), .ZN(_09694_ ) );
BUF_X4 _13242_ ( .A(_09611_ ), .Z(_09695_ ) );
NAND3_X1 _13243_ ( .A1(_09642_ ), .A2(_09136_ ), .A3(_09695_ ), .ZN(_09696_ ) );
AOI21_X1 _13244_ ( .A(fanout_net_8 ), .B1(_09694_ ), .B2(_09696_ ), .ZN(_00171_ ) );
OAI21_X1 _13245_ ( .A(\u_lsu.pmem[289] ), .B1(_09441_ ), .B2(_09648_ ), .ZN(_09697_ ) );
BUF_X4 _13246_ ( .A(_09616_ ), .Z(_09698_ ) );
NAND3_X1 _13247_ ( .A1(_09642_ ), .A2(_09136_ ), .A3(_09698_ ), .ZN(_09699_ ) );
AOI21_X1 _13248_ ( .A(fanout_net_8 ), .B1(_09697_ ), .B2(_09699_ ), .ZN(_00172_ ) );
INV_X4 _13249_ ( .A(_09145_ ), .ZN(_09700_ ) );
NAND3_X1 _13250_ ( .A1(_09700_ ), .A2(_08631_ ), .A3(_09125_ ), .ZN(_09701_ ) );
BUF_X4 _13251_ ( .A(_09535_ ), .Z(_09702_ ) );
NOR3_X4 _13252_ ( .A1(_09701_ ), .A2(_09702_ ), .A3(_09536_ ), .ZN(_09703_ ) );
NAND4_X1 _13253_ ( .A1(_09703_ ), .A2(_09672_ ), .A3(_09686_ ), .A4(_09676_ ), .ZN(_09704_ ) );
OAI21_X1 _13254_ ( .A(\u_lsu.pmem[288] ), .B1(_09441_ ), .B2(_09678_ ), .ZN(_09705_ ) );
AOI21_X1 _13255_ ( .A(fanout_net_9 ), .B1(_09704_ ), .B2(_09705_ ), .ZN(_00173_ ) );
BUF_X4 _13256_ ( .A(_09666_ ), .Z(_09706_ ) );
BUF_X2 _13257_ ( .A(_09465_ ), .Z(_09707_ ) );
AND3_X2 _13258_ ( .A1(_09566_ ), .A2(_09706_ ), .A3(_09707_ ), .ZN(_09708_ ) );
BUF_X4 _13259_ ( .A(_09675_ ), .Z(_09709_ ) );
NAND4_X1 _13260_ ( .A1(_09708_ ), .A2(_09672_ ), .A3(_09686_ ), .A4(_09709_ ), .ZN(_09710_ ) );
OAI21_X1 _13261_ ( .A(\u_lsu.pmem[263] ), .B1(_09469_ ), .B2(_09678_ ), .ZN(_09711_ ) );
AOI21_X1 _13262_ ( .A(fanout_net_9 ), .B1(_09710_ ), .B2(_09711_ ), .ZN(_00174_ ) );
OAI21_X1 _13263_ ( .A(\u_lsu.pmem[3973] ), .B1(_09599_ ), .B2(_09648_ ), .ZN(_09712_ ) );
BUF_X4 _13264_ ( .A(_09582_ ), .Z(_09713_ ) );
NAND4_X1 _13265_ ( .A1(_09602_ ), .A2(_09713_ ), .A3(_09659_ ), .A4(_09523_ ), .ZN(_09714_ ) );
AOI21_X1 _13266_ ( .A(fanout_net_9 ), .B1(_09712_ ), .B2(_09714_ ), .ZN(_00175_ ) );
AND3_X2 _13267_ ( .A1(_09578_ ), .A2(_09706_ ), .A3(_09707_ ), .ZN(_09715_ ) );
NAND4_X1 _13268_ ( .A1(_09715_ ), .A2(_09672_ ), .A3(_09686_ ), .A4(_09709_ ), .ZN(_09716_ ) );
OAI21_X1 _13269_ ( .A(\u_lsu.pmem[262] ), .B1(_09469_ ), .B2(_09678_ ), .ZN(_09717_ ) );
AOI21_X1 _13270_ ( .A(fanout_net_9 ), .B1(_09716_ ), .B2(_09717_ ), .ZN(_00176_ ) );
AND3_X2 _13271_ ( .A1(_09585_ ), .A2(_09706_ ), .A3(_09707_ ), .ZN(_09718_ ) );
NAND4_X1 _13272_ ( .A1(_09718_ ), .A2(_09672_ ), .A3(_09686_ ), .A4(_09709_ ), .ZN(_09719_ ) );
OAI21_X1 _13273_ ( .A(\u_lsu.pmem[261] ), .B1(_09469_ ), .B2(_09678_ ), .ZN(_09720_ ) );
AOI21_X1 _13274_ ( .A(fanout_net_9 ), .B1(_09719_ ), .B2(_09720_ ), .ZN(_00177_ ) );
AND3_X2 _13275_ ( .A1(_09148_ ), .A2(_09706_ ), .A3(_09707_ ), .ZN(_09721_ ) );
NAND4_X1 _13276_ ( .A1(_09721_ ), .A2(_09672_ ), .A3(_09686_ ), .A4(_09709_ ), .ZN(_09722_ ) );
OAI21_X1 _13277_ ( .A(\u_lsu.pmem[260] ), .B1(_09469_ ), .B2(_09678_ ), .ZN(_09723_ ) );
AOI21_X1 _13278_ ( .A(fanout_net_9 ), .B1(_09722_ ), .B2(_09723_ ), .ZN(_00178_ ) );
AND2_X1 _13279_ ( .A1(_09447_ ), .A2(_09465_ ), .ZN(_09724_ ) );
AND2_X2 _13280_ ( .A1(_09724_ ), .A2(_09667_ ), .ZN(_09725_ ) );
NAND4_X1 _13281_ ( .A1(_09725_ ), .A2(_09672_ ), .A3(_09686_ ), .A4(_09709_ ), .ZN(_09726_ ) );
OAI21_X1 _13282_ ( .A(\u_lsu.pmem[259] ), .B1(_09469_ ), .B2(_09678_ ), .ZN(_09727_ ) );
AOI21_X1 _13283_ ( .A(fanout_net_9 ), .B1(_09726_ ), .B2(_09727_ ), .ZN(_00179_ ) );
BUF_X4 _13284_ ( .A(_09459_ ), .Z(_09728_ ) );
NAND4_X1 _13285_ ( .A1(_09728_ ), .A2(_09474_ ), .A3(_09686_ ), .A4(_09467_ ), .ZN(_09729_ ) );
BUF_X8 _13286_ ( .A(_09450_ ), .Z(_09730_ ) );
BUF_X4 _13287_ ( .A(_09730_ ), .Z(_09731_ ) );
OAI21_X1 _13288_ ( .A(\u_lsu.pmem[258] ), .B1(_09469_ ), .B2(_09731_ ), .ZN(_09732_ ) );
AOI21_X1 _13289_ ( .A(fanout_net_9 ), .B1(_09729_ ), .B2(_09732_ ), .ZN(_00180_ ) );
AND3_X2 _13290_ ( .A1(_09616_ ), .A2(_09706_ ), .A3(_09707_ ), .ZN(_09733_ ) );
NAND4_X1 _13291_ ( .A1(_09733_ ), .A2(_09672_ ), .A3(_09686_ ), .A4(_09709_ ), .ZN(_09734_ ) );
OAI21_X1 _13292_ ( .A(\u_lsu.pmem[257] ), .B1(_09469_ ), .B2(_09731_ ), .ZN(_09735_ ) );
AOI21_X1 _13293_ ( .A(fanout_net_9 ), .B1(_09734_ ), .B2(_09735_ ), .ZN(_00181_ ) );
AND3_X2 _13294_ ( .A1(_09620_ ), .A2(_09706_ ), .A3(_09707_ ), .ZN(_09736_ ) );
BUF_X4 _13295_ ( .A(_09671_ ), .Z(_09737_ ) );
NAND4_X1 _13296_ ( .A1(_09736_ ), .A2(_09737_ ), .A3(_09686_ ), .A4(_09709_ ), .ZN(_09738_ ) );
OAI21_X1 _13297_ ( .A(\u_lsu.pmem[256] ), .B1(_09469_ ), .B2(_09731_ ), .ZN(_09739_ ) );
AOI21_X1 _13298_ ( .A(fanout_net_9 ), .B1(_09738_ ), .B2(_09739_ ), .ZN(_00182_ ) );
BUF_X4 _13299_ ( .A(_09456_ ), .Z(_09740_ ) );
BUF_X4 _13300_ ( .A(_09566_ ), .Z(_09741_ ) );
BUF_X4 _13301_ ( .A(_09741_ ), .Z(_09742_ ) );
BUF_X4 _13302_ ( .A(_09118_ ), .Z(_09743_ ) );
BUF_X4 _13303_ ( .A(_09550_ ), .Z(_09744_ ) );
BUF_X32 _13304_ ( .A(_09554_ ), .Z(_09745_ ) );
BUF_X4 _13305_ ( .A(_09745_ ), .Z(_09746_ ) );
AND2_X4 _13306_ ( .A1(_09084_ ), .A2(_09746_ ), .ZN(_09747_ ) );
NAND3_X1 _13307_ ( .A1(_09129_ ), .A2(_09744_ ), .A3(_09747_ ), .ZN(_09748_ ) );
NOR2_X1 _13308_ ( .A1(_09743_ ), .A2(_09748_ ), .ZN(_09749_ ) );
NAND4_X1 _13309_ ( .A1(_09728_ ), .A2(_09740_ ), .A3(_09742_ ), .A4(_09749_ ), .ZN(_09750_ ) );
NAND2_X1 _13310_ ( .A1(_09461_ ), .A2(_09749_ ), .ZN(_09751_ ) );
BUF_X4 _13311_ ( .A(_09751_ ), .Z(_09752_ ) );
OAI21_X1 _13312_ ( .A(\u_lsu.pmem[231] ), .B1(_09752_ ), .B2(_09731_ ), .ZN(_09753_ ) );
AOI21_X1 _13313_ ( .A(fanout_net_9 ), .B1(_09750_ ), .B2(_09753_ ), .ZN(_00183_ ) );
BUF_X2 _13314_ ( .A(_09747_ ), .Z(_09754_ ) );
AND3_X1 _13315_ ( .A1(_09577_ ), .A2(_09535_ ), .A3(_09754_ ), .ZN(_09755_ ) );
AND2_X2 _13316_ ( .A1(_09755_ ), .A2(_09667_ ), .ZN(_09756_ ) );
BUF_X4 _13317_ ( .A(_09673_ ), .Z(_09757_ ) );
NAND4_X1 _13318_ ( .A1(_09756_ ), .A2(_09737_ ), .A3(_09757_ ), .A4(_09709_ ), .ZN(_09758_ ) );
OAI21_X1 _13319_ ( .A(\u_lsu.pmem[230] ), .B1(_09752_ ), .B2(_09731_ ), .ZN(_09759_ ) );
AOI21_X1 _13320_ ( .A(fanout_net_9 ), .B1(_09758_ ), .B2(_09759_ ), .ZN(_00184_ ) );
BUF_X4 _13321_ ( .A(_09534_ ), .Z(_09760_ ) );
NAND3_X1 _13322_ ( .A1(_09585_ ), .A2(_09760_ ), .A3(_09754_ ), .ZN(_09761_ ) );
BUF_X4 _13323_ ( .A(_09536_ ), .Z(_09762_ ) );
NOR2_X1 _13324_ ( .A1(_09761_ ), .A2(_09762_ ), .ZN(_09763_ ) );
NAND4_X1 _13325_ ( .A1(_09763_ ), .A2(_09737_ ), .A3(_09757_ ), .A4(_09709_ ), .ZN(_09764_ ) );
OAI21_X1 _13326_ ( .A(\u_lsu.pmem[229] ), .B1(_09752_ ), .B2(_09731_ ), .ZN(_09765_ ) );
AOI21_X1 _13327_ ( .A(fanout_net_9 ), .B1(_09764_ ), .B2(_09765_ ), .ZN(_00185_ ) );
BUF_X4 _13328_ ( .A(_09647_ ), .Z(_09766_ ) );
OAI21_X1 _13329_ ( .A(\u_lsu.pmem[3972] ), .B1(_09599_ ), .B2(_09766_ ), .ZN(_09767_ ) );
NAND4_X1 _13330_ ( .A1(_09602_ ), .A2(_09514_ ), .A3(_09659_ ), .A4(_09523_ ), .ZN(_09768_ ) );
AOI21_X1 _13331_ ( .A(fanout_net_9 ), .B1(_09767_ ), .B2(_09768_ ), .ZN(_00186_ ) );
AND3_X1 _13332_ ( .A1(_09147_ ), .A2(_09535_ ), .A3(_09754_ ), .ZN(_09769_ ) );
AND2_X2 _13333_ ( .A1(_09769_ ), .A2(_09667_ ), .ZN(_09770_ ) );
NAND4_X1 _13334_ ( .A1(_09770_ ), .A2(_09737_ ), .A3(_09757_ ), .A4(_09709_ ), .ZN(_09771_ ) );
OAI21_X1 _13335_ ( .A(\u_lsu.pmem[228] ), .B1(_09752_ ), .B2(_09731_ ), .ZN(_09772_ ) );
AOI21_X1 _13336_ ( .A(fanout_net_9 ), .B1(_09771_ ), .B2(_09772_ ), .ZN(_00187_ ) );
NAND3_X1 _13337_ ( .A1(_09447_ ), .A2(_09760_ ), .A3(_09754_ ), .ZN(_09773_ ) );
BUF_X4 _13338_ ( .A(_09536_ ), .Z(_09774_ ) );
NOR2_X2 _13339_ ( .A1(_09773_ ), .A2(_09774_ ), .ZN(_09775_ ) );
BUF_X4 _13340_ ( .A(_09675_ ), .Z(_09776_ ) );
NAND4_X1 _13341_ ( .A1(_09775_ ), .A2(_09737_ ), .A3(_09757_ ), .A4(_09776_ ), .ZN(_09777_ ) );
OAI21_X1 _13342_ ( .A(\u_lsu.pmem[227] ), .B1(_09752_ ), .B2(_09731_ ), .ZN(_09778_ ) );
AOI21_X1 _13343_ ( .A(fanout_net_9 ), .B1(_09777_ ), .B2(_09778_ ), .ZN(_00188_ ) );
NAND3_X1 _13344_ ( .A1(_09610_ ), .A2(_09760_ ), .A3(_09754_ ), .ZN(_09779_ ) );
NOR2_X4 _13345_ ( .A1(_09779_ ), .A2(_09774_ ), .ZN(_09780_ ) );
NAND4_X1 _13346_ ( .A1(_09780_ ), .A2(_09737_ ), .A3(_09757_ ), .A4(_09776_ ), .ZN(_09781_ ) );
OAI21_X1 _13347_ ( .A(\u_lsu.pmem[226] ), .B1(_09752_ ), .B2(_09731_ ), .ZN(_09782_ ) );
AOI21_X1 _13348_ ( .A(fanout_net_9 ), .B1(_09781_ ), .B2(_09782_ ), .ZN(_00189_ ) );
NAND3_X1 _13349_ ( .A1(_09700_ ), .A2(_08638_ ), .A3(_09747_ ), .ZN(_09783_ ) );
BUF_X4 _13350_ ( .A(_09046_ ), .Z(_09784_ ) );
BUF_X4 _13351_ ( .A(_09784_ ), .Z(_09785_ ) );
BUF_X2 _13352_ ( .A(_09785_ ), .Z(\alu_result_out[6] ) );
BUF_X2 _13353_ ( .A(_09668_ ), .Z(_09786_ ) );
NOR3_X4 _13354_ ( .A1(_09783_ ), .A2(\alu_result_out[6] ), .A3(_09786_ ), .ZN(_09787_ ) );
NAND4_X1 _13355_ ( .A1(_09787_ ), .A2(_09737_ ), .A3(_09757_ ), .A4(_09776_ ), .ZN(_09788_ ) );
OAI21_X1 _13356_ ( .A(\u_lsu.pmem[225] ), .B1(_09752_ ), .B2(_09731_ ), .ZN(_09789_ ) );
AOI21_X1 _13357_ ( .A(fanout_net_9 ), .B1(_09788_ ), .B2(_09789_ ), .ZN(_00190_ ) );
NAND3_X1 _13358_ ( .A1(_09620_ ), .A2(_09760_ ), .A3(_09754_ ), .ZN(_09790_ ) );
NOR2_X2 _13359_ ( .A1(_09790_ ), .A2(_09774_ ), .ZN(_09791_ ) );
NAND4_X1 _13360_ ( .A1(_09791_ ), .A2(_09737_ ), .A3(_09757_ ), .A4(_09776_ ), .ZN(_09792_ ) );
BUF_X4 _13361_ ( .A(_09730_ ), .Z(_09793_ ) );
OAI21_X1 _13362_ ( .A(\u_lsu.pmem[224] ), .B1(_09752_ ), .B2(_09793_ ), .ZN(_09794_ ) );
AOI21_X1 _13363_ ( .A(fanout_net_9 ), .B1(_09792_ ), .B2(_09794_ ), .ZN(_00191_ ) );
BUF_X4 _13364_ ( .A(_09627_ ), .Z(_09795_ ) );
AND2_X4 _13365_ ( .A1(_09119_ ), .A2(_09795_ ), .ZN(_09796_ ) );
NAND3_X1 _13366_ ( .A1(_09129_ ), .A2(_09744_ ), .A3(_09796_ ), .ZN(_09797_ ) );
NOR2_X1 _13367_ ( .A1(_09743_ ), .A2(_09797_ ), .ZN(_09798_ ) );
NAND2_X1 _13368_ ( .A1(_09461_ ), .A2(_09798_ ), .ZN(_09799_ ) );
NOR2_X1 _13369_ ( .A1(_09799_ ), .A2(_09635_ ), .ZN(_09800_ ) );
OAI21_X1 _13370_ ( .A(_09110_ ), .B1(_09800_ ), .B2(\u_lsu.pmem[199] ), .ZN(_09801_ ) );
AOI21_X1 _13371_ ( .A(_09801_ ), .B1(_09638_ ), .B2(_09800_ ), .ZN(_00192_ ) );
CLKBUF_X2 _13372_ ( .A(_09796_ ), .Z(_09802_ ) );
NAND3_X1 _13373_ ( .A1(_09578_ ), .A2(_09702_ ), .A3(_09802_ ), .ZN(_09803_ ) );
NOR2_X4 _13374_ ( .A1(_09803_ ), .A2(\alu_result_out[6] ), .ZN(_09804_ ) );
BUF_X4 _13375_ ( .A(_08995_ ), .Z(_09805_ ) );
BUF_X4 _13376_ ( .A(_09805_ ), .Z(_09806_ ) );
NAND4_X1 _13377_ ( .A1(_09804_ ), .A2(_09806_ ), .A3(_09757_ ), .A4(_09776_ ), .ZN(_09807_ ) );
BUF_X4 _13378_ ( .A(_09799_ ), .Z(_09808_ ) );
OAI21_X1 _13379_ ( .A(\u_lsu.pmem[198] ), .B1(_09808_ ), .B2(_09793_ ), .ZN(_09809_ ) );
AOI21_X1 _13380_ ( .A(fanout_net_9 ), .B1(_09807_ ), .B2(_09809_ ), .ZN(_00193_ ) );
NAND3_X1 _13381_ ( .A1(_09584_ ), .A2(_09702_ ), .A3(_09802_ ), .ZN(_09810_ ) );
NOR2_X1 _13382_ ( .A1(_09810_ ), .A2(_09774_ ), .ZN(_09811_ ) );
NAND4_X1 _13383_ ( .A1(_09811_ ), .A2(_09737_ ), .A3(_09757_ ), .A4(_09776_ ), .ZN(_09812_ ) );
OAI21_X1 _13384_ ( .A(\u_lsu.pmem[197] ), .B1(_09808_ ), .B2(_09793_ ), .ZN(_09813_ ) );
AOI21_X1 _13385_ ( .A(fanout_net_9 ), .B1(_09812_ ), .B2(_09813_ ), .ZN(_00194_ ) );
AND3_X1 _13386_ ( .A1(_09147_ ), .A2(_09535_ ), .A3(_09802_ ), .ZN(_09814_ ) );
AND2_X2 _13387_ ( .A1(_09814_ ), .A2(_09667_ ), .ZN(_09815_ ) );
NAND4_X1 _13388_ ( .A1(_09815_ ), .A2(_09737_ ), .A3(_09757_ ), .A4(_09776_ ), .ZN(_09816_ ) );
OAI21_X1 _13389_ ( .A(\u_lsu.pmem[196] ), .B1(_09808_ ), .B2(_09793_ ), .ZN(_09817_ ) );
AOI21_X1 _13390_ ( .A(fanout_net_9 ), .B1(_09816_ ), .B2(_09817_ ), .ZN(_00195_ ) );
AND3_X1 _13391_ ( .A1(_09447_ ), .A2(_09535_ ), .A3(_09802_ ), .ZN(_09818_ ) );
AND2_X2 _13392_ ( .A1(_09818_ ), .A2(_09667_ ), .ZN(_09819_ ) );
BUF_X4 _13393_ ( .A(_09671_ ), .Z(_09820_ ) );
BUF_X4 _13394_ ( .A(_09673_ ), .Z(_09821_ ) );
NAND4_X1 _13395_ ( .A1(_09819_ ), .A2(_09820_ ), .A3(_09821_ ), .A4(_09776_ ), .ZN(_09822_ ) );
OAI21_X1 _13396_ ( .A(\u_lsu.pmem[195] ), .B1(_09808_ ), .B2(_09793_ ), .ZN(_09823_ ) );
AOI21_X1 _13397_ ( .A(fanout_net_9 ), .B1(_09822_ ), .B2(_09823_ ), .ZN(_00196_ ) );
OAI21_X1 _13398_ ( .A(\u_lsu.pmem[3971] ), .B1(_09599_ ), .B2(_09766_ ), .ZN(_09824_ ) );
NAND4_X1 _13399_ ( .A1(_09602_ ), .A2(_09520_ ), .A3(_09659_ ), .A4(_09523_ ), .ZN(_09825_ ) );
AOI21_X1 _13400_ ( .A(fanout_net_9 ), .B1(_09824_ ), .B2(_09825_ ), .ZN(_00197_ ) );
NAND3_X1 _13401_ ( .A1(_09610_ ), .A2(_09702_ ), .A3(_09802_ ), .ZN(_09826_ ) );
NOR2_X4 _13402_ ( .A1(_09826_ ), .A2(_09774_ ), .ZN(_09827_ ) );
NAND4_X1 _13403_ ( .A1(_09827_ ), .A2(_09820_ ), .A3(_09821_ ), .A4(_09776_ ), .ZN(_09828_ ) );
OAI21_X1 _13404_ ( .A(\u_lsu.pmem[194] ), .B1(_09808_ ), .B2(_09793_ ), .ZN(_09829_ ) );
AOI21_X1 _13405_ ( .A(fanout_net_9 ), .B1(_09828_ ), .B2(_09829_ ), .ZN(_00198_ ) );
NAND3_X1 _13406_ ( .A1(_09700_ ), .A2(_08638_ ), .A3(_09796_ ), .ZN(_09830_ ) );
NOR3_X4 _13407_ ( .A1(_09830_ ), .A2(_09785_ ), .A3(_09786_ ), .ZN(_09831_ ) );
NAND4_X1 _13408_ ( .A1(_09831_ ), .A2(_09820_ ), .A3(_09821_ ), .A4(_09776_ ), .ZN(_09832_ ) );
OAI21_X1 _13409_ ( .A(\u_lsu.pmem[193] ), .B1(_09808_ ), .B2(_09793_ ), .ZN(_09833_ ) );
AOI21_X1 _13410_ ( .A(fanout_net_9 ), .B1(_09832_ ), .B2(_09833_ ), .ZN(_00199_ ) );
NAND3_X1 _13411_ ( .A1(_09620_ ), .A2(_09702_ ), .A3(_09802_ ), .ZN(_09834_ ) );
NOR2_X2 _13412_ ( .A1(_09834_ ), .A2(_09774_ ), .ZN(_09835_ ) );
BUF_X4 _13413_ ( .A(_09675_ ), .Z(_09836_ ) );
NAND4_X1 _13414_ ( .A1(_09835_ ), .A2(_09820_ ), .A3(_09821_ ), .A4(_09836_ ), .ZN(_09837_ ) );
OAI21_X1 _13415_ ( .A(\u_lsu.pmem[192] ), .B1(_09808_ ), .B2(_09793_ ), .ZN(_09838_ ) );
AOI21_X1 _13416_ ( .A(fanout_net_9 ), .B1(_09837_ ), .B2(_09838_ ), .ZN(_00200_ ) );
NAND3_X1 _13417_ ( .A1(_09566_ ), .A2(_09702_ ), .A3(_09485_ ), .ZN(_09839_ ) );
NOR2_X1 _13418_ ( .A1(_09839_ ), .A2(_09774_ ), .ZN(_09840_ ) );
NAND4_X1 _13419_ ( .A1(_09840_ ), .A2(_09820_ ), .A3(_09821_ ), .A4(_09836_ ), .ZN(_09841_ ) );
BUF_X4 _13420_ ( .A(_09506_ ), .Z(_09842_ ) );
AND2_X1 _13421_ ( .A1(_09463_ ), .A2(_09485_ ), .ZN(_09843_ ) );
AND2_X1 _13422_ ( .A1(_09505_ ), .A2(_09843_ ), .ZN(_09844_ ) );
NAND3_X1 _13423_ ( .A1(_09454_ ), .A2(_09842_ ), .A3(_09844_ ), .ZN(_09845_ ) );
BUF_X4 _13424_ ( .A(_09845_ ), .Z(_09846_ ) );
OAI21_X1 _13425_ ( .A(\u_lsu.pmem[167] ), .B1(_09846_ ), .B2(_09793_ ), .ZN(_09847_ ) );
AOI21_X1 _13426_ ( .A(fanout_net_9 ), .B1(_09841_ ), .B2(_09847_ ), .ZN(_00201_ ) );
NAND3_X1 _13427_ ( .A1(_09577_ ), .A2(_09702_ ), .A3(_09485_ ), .ZN(_09848_ ) );
NOR2_X1 _13428_ ( .A1(_09848_ ), .A2(_09774_ ), .ZN(_09849_ ) );
NAND4_X1 _13429_ ( .A1(_09849_ ), .A2(_09820_ ), .A3(_09821_ ), .A4(_09836_ ), .ZN(_09850_ ) );
OAI21_X1 _13430_ ( .A(\u_lsu.pmem[166] ), .B1(_09846_ ), .B2(_09793_ ), .ZN(_09851_ ) );
AOI21_X1 _13431_ ( .A(fanout_net_9 ), .B1(_09850_ ), .B2(_09851_ ), .ZN(_00202_ ) );
NAND3_X1 _13432_ ( .A1(_09584_ ), .A2(_09702_ ), .A3(_09485_ ), .ZN(_09852_ ) );
NOR2_X1 _13433_ ( .A1(_09852_ ), .A2(_09774_ ), .ZN(_09853_ ) );
NAND4_X1 _13434_ ( .A1(_09853_ ), .A2(_09820_ ), .A3(_09821_ ), .A4(_09836_ ), .ZN(_09854_ ) );
BUF_X4 _13435_ ( .A(_09730_ ), .Z(_09855_ ) );
OAI21_X1 _13436_ ( .A(\u_lsu.pmem[165] ), .B1(_09846_ ), .B2(_09855_ ), .ZN(_09856_ ) );
AOI21_X1 _13437_ ( .A(fanout_net_9 ), .B1(_09854_ ), .B2(_09856_ ), .ZN(_00203_ ) );
BUF_X4 _13438_ ( .A(_09843_ ), .Z(_09857_ ) );
AND3_X2 _13439_ ( .A1(_09148_ ), .A2(_09706_ ), .A3(_09857_ ), .ZN(_09858_ ) );
NAND4_X1 _13440_ ( .A1(_09858_ ), .A2(_09820_ ), .A3(_09821_ ), .A4(_09836_ ), .ZN(_09859_ ) );
OAI21_X1 _13441_ ( .A(\u_lsu.pmem[164] ), .B1(_09846_ ), .B2(_09855_ ), .ZN(_09860_ ) );
AOI21_X1 _13442_ ( .A(fanout_net_10 ), .B1(_09859_ ), .B2(_09860_ ), .ZN(_00204_ ) );
AND3_X2 _13443_ ( .A1(_09447_ ), .A2(_09706_ ), .A3(_09857_ ), .ZN(_09861_ ) );
NAND4_X1 _13444_ ( .A1(_09861_ ), .A2(_09820_ ), .A3(_09821_ ), .A4(_09836_ ), .ZN(_09862_ ) );
OAI21_X1 _13445_ ( .A(\u_lsu.pmem[163] ), .B1(_09846_ ), .B2(_09855_ ), .ZN(_09863_ ) );
AOI21_X1 _13446_ ( .A(fanout_net_10 ), .B1(_09862_ ), .B2(_09863_ ), .ZN(_00205_ ) );
AND3_X2 _13447_ ( .A1(_09611_ ), .A2(_09706_ ), .A3(_09857_ ), .ZN(_09864_ ) );
NAND4_X1 _13448_ ( .A1(_09864_ ), .A2(_09820_ ), .A3(_09821_ ), .A4(_09836_ ), .ZN(_09865_ ) );
OAI21_X1 _13449_ ( .A(\u_lsu.pmem[162] ), .B1(_09846_ ), .B2(_09855_ ), .ZN(_09866_ ) );
AOI21_X1 _13450_ ( .A(fanout_net_10 ), .B1(_09865_ ), .B2(_09866_ ), .ZN(_00206_ ) );
AND3_X2 _13451_ ( .A1(_09615_ ), .A2(_09706_ ), .A3(_09857_ ), .ZN(_09867_ ) );
BUF_X4 _13452_ ( .A(_09671_ ), .Z(_09868_ ) );
BUF_X4 _13453_ ( .A(_09673_ ), .Z(_09869_ ) );
NAND4_X1 _13454_ ( .A1(_09867_ ), .A2(_09868_ ), .A3(_09869_ ), .A4(_09836_ ), .ZN(_09870_ ) );
OAI21_X1 _13455_ ( .A(\u_lsu.pmem[161] ), .B1(_09846_ ), .B2(_09855_ ), .ZN(_09871_ ) );
AOI21_X1 _13456_ ( .A(fanout_net_10 ), .B1(_09870_ ), .B2(_09871_ ), .ZN(_00207_ ) );
OAI21_X1 _13457_ ( .A(\u_lsu.pmem[3970] ), .B1(_09599_ ), .B2(_09766_ ), .ZN(_09872_ ) );
BUF_X4 _13458_ ( .A(_09505_ ), .Z(_09873_ ) );
NOR3_X1 _13459_ ( .A1(_09533_ ), .A2(_09535_ ), .A3(_09873_ ), .ZN(_09874_ ) );
BUF_X8 _13460_ ( .A(_09743_ ), .Z(_09875_ ) );
BUF_X4 _13461_ ( .A(_09875_ ), .Z(_09876_ ) );
BUF_X8 _13462_ ( .A(_09135_ ), .Z(_09877_ ) );
BUF_X8 _13463_ ( .A(_09877_ ), .Z(_09878_ ) );
BUF_X4 _13464_ ( .A(_09878_ ), .Z(_09879_ ) );
NAND4_X1 _13465_ ( .A1(_09874_ ), .A2(_09876_ ), .A3(_09879_ ), .A4(_09523_ ), .ZN(_09880_ ) );
AOI21_X1 _13466_ ( .A(fanout_net_10 ), .B1(_09872_ ), .B2(_09880_ ), .ZN(_00208_ ) );
AND2_X2 _13467_ ( .A1(_09620_ ), .A2(_09844_ ), .ZN(_09881_ ) );
BUF_X4 _13468_ ( .A(_09675_ ), .Z(_09882_ ) );
BUF_X8 _13469_ ( .A(_09539_ ), .Z(_09883_ ) );
BUF_X4 _13470_ ( .A(_09883_ ), .Z(_09884_ ) );
BUF_X4 _13471_ ( .A(_09476_ ), .Z(_09885_ ) );
NAND4_X1 _13472_ ( .A1(_09881_ ), .A2(_09882_ ), .A3(_09884_ ), .A4(_09885_ ), .ZN(_09886_ ) );
OAI21_X1 _13473_ ( .A(\u_lsu.pmem[160] ), .B1(_09846_ ), .B2(_09855_ ), .ZN(_09887_ ) );
AOI21_X1 _13474_ ( .A(fanout_net_10 ), .B1(_09886_ ), .B2(_09887_ ), .ZN(_00209_ ) );
BUF_X4 _13475_ ( .A(_09744_ ), .Z(_09888_ ) );
NAND3_X4 _13476_ ( .A1(_09503_ ), .A2(_09888_ ), .A3(_09505_ ), .ZN(_09889_ ) );
OR3_X2 _13477_ ( .A1(_09889_ ), .A2(_09743_ ), .A3(_09135_ ), .ZN(_09890_ ) );
BUF_X4 _13478_ ( .A(_09890_ ), .Z(_09891_ ) );
OAI21_X1 _13479_ ( .A(\u_lsu.pmem[135] ), .B1(_09891_ ), .B2(_09766_ ), .ZN(_09892_ ) );
NOR2_X2 _13480_ ( .A1(_09889_ ), .A2(_09875_ ), .ZN(_09893_ ) );
BUF_X4 _13481_ ( .A(_09893_ ), .Z(_09894_ ) );
BUF_X4 _13482_ ( .A(_09522_ ), .Z(_09895_ ) );
NAND4_X1 _13483_ ( .A1(_09894_ ), .A2(_09603_ ), .A3(_09521_ ), .A4(_09895_ ), .ZN(_09896_ ) );
AOI21_X1 _13484_ ( .A(fanout_net_10 ), .B1(_09892_ ), .B2(_09896_ ), .ZN(_00210_ ) );
OAI21_X1 _13485_ ( .A(\u_lsu.pmem[134] ), .B1(_09891_ ), .B2(_09766_ ), .ZN(_09897_ ) );
NAND4_X1 _13486_ ( .A1(_09894_ ), .A2(_09658_ ), .A3(_09521_ ), .A4(_09895_ ), .ZN(_09898_ ) );
AOI21_X1 _13487_ ( .A(fanout_net_10 ), .B1(_09897_ ), .B2(_09898_ ), .ZN(_00211_ ) );
OAI21_X1 _13488_ ( .A(\u_lsu.pmem[133] ), .B1(_09891_ ), .B2(_09766_ ), .ZN(_09899_ ) );
NAND4_X1 _13489_ ( .A1(_09894_ ), .A2(_09713_ ), .A3(_09521_ ), .A4(_09895_ ), .ZN(_09900_ ) );
AOI21_X1 _13490_ ( .A(fanout_net_10 ), .B1(_09899_ ), .B2(_09900_ ), .ZN(_00212_ ) );
OAI21_X1 _13491_ ( .A(\u_lsu.pmem[132] ), .B1(_09891_ ), .B2(_09766_ ), .ZN(_09901_ ) );
NAND4_X1 _13492_ ( .A1(_09894_ ), .A2(_09514_ ), .A3(_09521_ ), .A4(_09895_ ), .ZN(_09902_ ) );
AOI21_X1 _13493_ ( .A(fanout_net_10 ), .B1(_09901_ ), .B2(_09902_ ), .ZN(_00213_ ) );
OAI21_X1 _13494_ ( .A(\u_lsu.pmem[131] ), .B1(_09891_ ), .B2(_09766_ ), .ZN(_09903_ ) );
NAND4_X1 _13495_ ( .A1(_09894_ ), .A2(_09520_ ), .A3(_09521_ ), .A4(_09895_ ), .ZN(_09904_ ) );
AOI21_X1 _13496_ ( .A(fanout_net_10 ), .B1(_09903_ ), .B2(_09904_ ), .ZN(_00214_ ) );
OAI21_X1 _13497_ ( .A(\u_lsu.pmem[130] ), .B1(_09891_ ), .B2(_09766_ ), .ZN(_09905_ ) );
NOR3_X1 _13498_ ( .A1(_09533_ ), .A2(_09785_ ), .A3(_09786_ ), .ZN(_09906_ ) );
NAND4_X1 _13499_ ( .A1(_09906_ ), .A2(_09540_ ), .A3(_09521_ ), .A4(_09895_ ), .ZN(_09907_ ) );
AOI21_X1 _13500_ ( .A(fanout_net_10 ), .B1(_09905_ ), .B2(_09907_ ), .ZN(_00215_ ) );
OAI21_X1 _13501_ ( .A(\u_lsu.pmem[129] ), .B1(_09891_ ), .B2(_09766_ ), .ZN(_09908_ ) );
BUF_X4 _13502_ ( .A(_09476_ ), .Z(_09909_ ) );
NAND4_X1 _13503_ ( .A1(_09894_ ), .A2(_09544_ ), .A3(_09909_ ), .A4(_09895_ ), .ZN(_09910_ ) );
AOI21_X1 _13504_ ( .A(fanout_net_10 ), .B1(_09908_ ), .B2(_09910_ ), .ZN(_00216_ ) );
BUF_X4 _13505_ ( .A(_09647_ ), .Z(_09911_ ) );
OAI21_X1 _13506_ ( .A(\u_lsu.pmem[128] ), .B1(_09891_ ), .B2(_09911_ ), .ZN(_09912_ ) );
NAND4_X1 _13507_ ( .A1(_09894_ ), .A2(_09548_ ), .A3(_09909_ ), .A4(_09895_ ), .ZN(_09913_ ) );
AOI21_X1 _13508_ ( .A(fanout_net_10 ), .B1(_09912_ ), .B2(_09913_ ), .ZN(_00217_ ) );
BUF_X4 _13509_ ( .A(_09566_ ), .Z(_09914_ ) );
AND3_X1 _13510_ ( .A1(_09129_ ), .A2(_09534_ ), .A3(_09556_ ), .ZN(_09915_ ) );
AND2_X2 _13511_ ( .A1(_09538_ ), .A2(_09915_ ), .ZN(_09916_ ) );
BUF_X4 _13512_ ( .A(_09916_ ), .Z(_09917_ ) );
NAND4_X1 _13513_ ( .A1(_09728_ ), .A2(_09740_ ), .A3(_09914_ ), .A4(_09917_ ), .ZN(_09918_ ) );
NAND2_X1 _13514_ ( .A1(_09916_ ), .A2(_09475_ ), .ZN(_09919_ ) );
BUF_X4 _13515_ ( .A(_09919_ ), .Z(_09920_ ) );
OAI21_X1 _13516_ ( .A(\u_lsu.pmem[103] ), .B1(_09920_ ), .B2(_09855_ ), .ZN(_09921_ ) );
AOI21_X1 _13517_ ( .A(fanout_net_10 ), .B1(_09918_ ), .B2(_09921_ ), .ZN(_00218_ ) );
OAI21_X1 _13518_ ( .A(\u_lsu.pmem[3969] ), .B1(_09599_ ), .B2(_09911_ ), .ZN(_09922_ ) );
BUF_X4 _13519_ ( .A(_09543_ ), .Z(_09923_ ) );
NAND4_X1 _13520_ ( .A1(_09602_ ), .A2(_09923_ ), .A3(_09659_ ), .A4(_09895_ ), .ZN(_09924_ ) );
AOI21_X1 _13521_ ( .A(fanout_net_10 ), .B1(_09922_ ), .B2(_09924_ ), .ZN(_00219_ ) );
BUF_X4 _13522_ ( .A(_09578_ ), .Z(_09925_ ) );
NAND4_X1 _13523_ ( .A1(_09728_ ), .A2(_09740_ ), .A3(_09925_ ), .A4(_09917_ ), .ZN(_09926_ ) );
OAI21_X1 _13524_ ( .A(\u_lsu.pmem[102] ), .B1(_09920_ ), .B2(_09855_ ), .ZN(_09927_ ) );
AOI21_X1 _13525_ ( .A(fanout_net_10 ), .B1(_09926_ ), .B2(_09927_ ), .ZN(_00220_ ) );
BUF_X4 _13526_ ( .A(_09585_ ), .Z(_09928_ ) );
NAND4_X1 _13527_ ( .A1(_09728_ ), .A2(_09740_ ), .A3(_09928_ ), .A4(_09917_ ), .ZN(_09929_ ) );
OAI21_X1 _13528_ ( .A(\u_lsu.pmem[101] ), .B1(_09920_ ), .B2(_09855_ ), .ZN(_09930_ ) );
AOI21_X1 _13529_ ( .A(fanout_net_10 ), .B1(_09929_ ), .B2(_09930_ ), .ZN(_00221_ ) );
BUF_X4 _13530_ ( .A(_09148_ ), .Z(_09931_ ) );
NAND4_X1 _13531_ ( .A1(_09728_ ), .A2(_09740_ ), .A3(_09931_ ), .A4(_09917_ ), .ZN(_09932_ ) );
OAI21_X1 _13532_ ( .A(\u_lsu.pmem[100] ), .B1(_09920_ ), .B2(_09855_ ), .ZN(_09933_ ) );
AOI21_X1 _13533_ ( .A(fanout_net_10 ), .B1(_09932_ ), .B2(_09933_ ), .ZN(_00222_ ) );
BUF_X4 _13534_ ( .A(_09448_ ), .Z(_09934_ ) );
NAND4_X1 _13535_ ( .A1(_09728_ ), .A2(_09740_ ), .A3(_09934_ ), .A4(_09917_ ), .ZN(_09935_ ) );
BUF_X4 _13536_ ( .A(_09730_ ), .Z(_09936_ ) );
OAI21_X1 _13537_ ( .A(\u_lsu.pmem[99] ), .B1(_09920_ ), .B2(_09936_ ), .ZN(_09937_ ) );
AOI21_X1 _13538_ ( .A(fanout_net_10 ), .B1(_09935_ ), .B2(_09937_ ), .ZN(_00223_ ) );
BUF_X4 _13539_ ( .A(_09611_ ), .Z(_09938_ ) );
NAND4_X1 _13540_ ( .A1(_09728_ ), .A2(_09740_ ), .A3(_09938_ ), .A4(_09917_ ), .ZN(_09939_ ) );
OAI21_X1 _13541_ ( .A(\u_lsu.pmem[98] ), .B1(_09920_ ), .B2(_09936_ ), .ZN(_09940_ ) );
AOI21_X1 _13542_ ( .A(fanout_net_10 ), .B1(_09939_ ), .B2(_09940_ ), .ZN(_00224_ ) );
BUF_X4 _13543_ ( .A(_09616_ ), .Z(_09941_ ) );
NAND4_X1 _13544_ ( .A1(_09728_ ), .A2(_09740_ ), .A3(_09941_ ), .A4(_09917_ ), .ZN(_09942_ ) );
OAI21_X1 _13545_ ( .A(\u_lsu.pmem[97] ), .B1(_09920_ ), .B2(_09936_ ), .ZN(_09943_ ) );
AOI21_X1 _13546_ ( .A(fanout_net_10 ), .B1(_09942_ ), .B2(_09943_ ), .ZN(_00225_ ) );
BUF_X4 _13547_ ( .A(_09621_ ), .Z(_09944_ ) );
NAND4_X1 _13548_ ( .A1(_09728_ ), .A2(_09740_ ), .A3(_09944_ ), .A4(_09917_ ), .ZN(_09945_ ) );
OAI21_X1 _13549_ ( .A(\u_lsu.pmem[96] ), .B1(_09920_ ), .B2(_09936_ ), .ZN(_09946_ ) );
AOI21_X1 _13550_ ( .A(fanout_net_10 ), .B1(_09945_ ), .B2(_09946_ ), .ZN(_00226_ ) );
AND2_X1 _13551_ ( .A1(_09055_ ), .A2(_09629_ ), .ZN(_09947_ ) );
AND2_X4 _13552_ ( .A1(_09129_ ), .A2(_09947_ ), .ZN(_09948_ ) );
NAND3_X4 _13553_ ( .A1(_09454_ ), .A2(_09842_ ), .A3(_09948_ ), .ZN(_09949_ ) );
BUF_X4 _13554_ ( .A(_09140_ ), .Z(_09950_ ) );
NOR2_X1 _13555_ ( .A1(_09949_ ), .A2(_09950_ ), .ZN(_09951_ ) );
NOR2_X1 _13556_ ( .A1(_09951_ ), .A2(\u_lsu.pmem[71] ), .ZN(_09952_ ) );
AOI211_X1 _13557_ ( .A(fanout_net_10 ), .B(_09952_ ), .C1(_09568_ ), .C2(_09951_ ), .ZN(_00227_ ) );
BUF_X8 _13558_ ( .A(_09458_ ), .Z(_09953_ ) );
BUF_X4 _13559_ ( .A(_09953_ ), .Z(_09954_ ) );
BUF_X4 _13560_ ( .A(_09145_ ), .Z(_09955_ ) );
INV_X1 _13561_ ( .A(_09948_ ), .ZN(_09956_ ) );
NOR3_X2 _13562_ ( .A1(_09955_ ), .A2(_09576_ ), .A3(_09956_ ), .ZN(_09957_ ) );
NAND4_X1 _13563_ ( .A1(_09954_ ), .A2(_09957_ ), .A3(_09884_ ), .A4(_09885_ ), .ZN(_09958_ ) );
BUF_X4 _13564_ ( .A(_09949_ ), .Z(_09959_ ) );
OAI21_X1 _13565_ ( .A(\u_lsu.pmem[70] ), .B1(_09959_ ), .B2(_09936_ ), .ZN(_09960_ ) );
AOI21_X1 _13566_ ( .A(fanout_net_10 ), .B1(_09958_ ), .B2(_09960_ ), .ZN(_00228_ ) );
NOR3_X2 _13567_ ( .A1(_09955_ ), .A2(_09583_ ), .A3(_09956_ ), .ZN(_09961_ ) );
NAND4_X1 _13568_ ( .A1(_09954_ ), .A2(_09961_ ), .A3(_09884_ ), .A4(_09885_ ), .ZN(_09962_ ) );
OAI21_X1 _13569_ ( .A(\u_lsu.pmem[69] ), .B1(_09959_ ), .B2(_09936_ ), .ZN(_09963_ ) );
AOI21_X1 _13570_ ( .A(fanout_net_10 ), .B1(_09962_ ), .B2(_09963_ ), .ZN(_00229_ ) );
OAI21_X1 _13571_ ( .A(\u_lsu.pmem[3968] ), .B1(_09599_ ), .B2(_09911_ ), .ZN(_09964_ ) );
NAND4_X1 _13572_ ( .A1(_09601_ ), .A2(_09548_ ), .A3(_09659_ ), .A4(_09895_ ), .ZN(_09965_ ) );
AOI21_X1 _13573_ ( .A(fanout_net_10 ), .B1(_09964_ ), .B2(_09965_ ), .ZN(_00230_ ) );
NOR3_X2 _13574_ ( .A1(_09955_ ), .A2(_09146_ ), .A3(_09956_ ), .ZN(_09966_ ) );
NAND4_X1 _13575_ ( .A1(_09954_ ), .A2(_09966_ ), .A3(_09884_ ), .A4(_09885_ ), .ZN(_09967_ ) );
OAI21_X1 _13576_ ( .A(\u_lsu.pmem[68] ), .B1(_09959_ ), .B2(_09936_ ), .ZN(_09968_ ) );
AOI21_X1 _13577_ ( .A(fanout_net_10 ), .B1(_09967_ ), .B2(_09968_ ), .ZN(_00231_ ) );
CLKBUF_X2 _13578_ ( .A(_09446_ ), .Z(_09969_ ) );
NOR3_X2 _13579_ ( .A1(_09955_ ), .A2(_09969_ ), .A3(_09956_ ), .ZN(_09970_ ) );
NAND4_X1 _13580_ ( .A1(_09954_ ), .A2(_09970_ ), .A3(_09884_ ), .A4(_09885_ ), .ZN(_09971_ ) );
OAI21_X1 _13581_ ( .A(\u_lsu.pmem[67] ), .B1(_09959_ ), .B2(_09936_ ), .ZN(_09972_ ) );
AOI21_X1 _13582_ ( .A(fanout_net_10 ), .B1(_09971_ ), .B2(_09972_ ), .ZN(_00232_ ) );
CLKBUF_X2 _13583_ ( .A(_08962_ ), .Z(_09973_ ) );
NOR3_X2 _13584_ ( .A1(_09145_ ), .A2(_09973_ ), .A3(_09956_ ), .ZN(_09974_ ) );
NAND4_X1 _13585_ ( .A1(_09954_ ), .A2(_09974_ ), .A3(_09884_ ), .A4(_09885_ ), .ZN(_09975_ ) );
OAI21_X1 _13586_ ( .A(\u_lsu.pmem[66] ), .B1(_09959_ ), .B2(_09936_ ), .ZN(_09976_ ) );
AOI21_X1 _13587_ ( .A(fanout_net_10 ), .B1(_09975_ ), .B2(_09976_ ), .ZN(_00233_ ) );
CLKBUF_X2 _13588_ ( .A(_08639_ ), .Z(_09977_ ) );
NOR3_X2 _13589_ ( .A1(_09145_ ), .A2(_09977_ ), .A3(_09956_ ), .ZN(_09978_ ) );
BUF_X4 _13590_ ( .A(_09883_ ), .Z(_09979_ ) );
NAND4_X1 _13591_ ( .A1(_09954_ ), .A2(_09978_ ), .A3(_09979_ ), .A4(_09885_ ), .ZN(_09980_ ) );
OAI21_X1 _13592_ ( .A(\u_lsu.pmem[65] ), .B1(_09959_ ), .B2(_09936_ ), .ZN(_09981_ ) );
AOI21_X1 _13593_ ( .A(fanout_net_11 ), .B1(_09980_ ), .B2(_09981_ ), .ZN(_00234_ ) );
NOR3_X2 _13594_ ( .A1(_09145_ ), .A2(_08952_ ), .A3(_09956_ ), .ZN(_09982_ ) );
NAND4_X1 _13595_ ( .A1(_09954_ ), .A2(_09982_ ), .A3(_09979_ ), .A4(_09885_ ), .ZN(_09983_ ) );
BUF_X4 _13596_ ( .A(_09730_ ), .Z(_09984_ ) );
OAI21_X1 _13597_ ( .A(\u_lsu.pmem[64] ), .B1(_09959_ ), .B2(_09984_ ), .ZN(_09985_ ) );
AOI21_X1 _13598_ ( .A(fanout_net_11 ), .B1(_09983_ ), .B2(_09985_ ), .ZN(_00235_ ) );
BUF_X4 _13599_ ( .A(_09873_ ), .Z(_09986_ ) );
AND3_X2 _13600_ ( .A1(_09663_ ), .A2(_09760_ ), .A3(_09986_ ), .ZN(_09987_ ) );
NAND4_X1 _13601_ ( .A1(_09987_ ), .A2(_09868_ ), .A3(_09869_ ), .A4(_09836_ ), .ZN(_09988_ ) );
AND3_X1 _13602_ ( .A1(_09129_ ), .A2(_09125_ ), .A3(_09534_ ), .ZN(_09989_ ) );
AND2_X1 _13603_ ( .A1(_09538_ ), .A2(_09989_ ), .ZN(_09990_ ) );
NAND2_X1 _13604_ ( .A1(_09990_ ), .A2(_09475_ ), .ZN(_09991_ ) );
BUF_X4 _13605_ ( .A(_09991_ ), .Z(_09992_ ) );
OAI21_X1 _13606_ ( .A(\u_lsu.pmem[39] ), .B1(_09992_ ), .B2(_09984_ ), .ZN(_09993_ ) );
AOI21_X1 _13607_ ( .A(fanout_net_11 ), .B1(_09988_ ), .B2(_09993_ ), .ZN(_00236_ ) );
AND3_X2 _13608_ ( .A1(_09680_ ), .A2(_09760_ ), .A3(_09986_ ), .ZN(_09994_ ) );
NAND4_X1 _13609_ ( .A1(_09994_ ), .A2(_09868_ ), .A3(_09869_ ), .A4(_09836_ ), .ZN(_09995_ ) );
OAI21_X1 _13610_ ( .A(\u_lsu.pmem[38] ), .B1(_09992_ ), .B2(_09984_ ), .ZN(_09996_ ) );
AOI21_X1 _13611_ ( .A(fanout_net_11 ), .B1(_09995_ ), .B2(_09996_ ), .ZN(_00237_ ) );
AND3_X2 _13612_ ( .A1(_09684_ ), .A2(_09760_ ), .A3(_09986_ ), .ZN(_09997_ ) );
BUF_X4 _13613_ ( .A(_09675_ ), .Z(_09998_ ) );
NAND4_X1 _13614_ ( .A1(_09997_ ), .A2(_09868_ ), .A3(_09869_ ), .A4(_09998_ ), .ZN(_09999_ ) );
OAI21_X1 _13615_ ( .A(\u_lsu.pmem[37] ), .B1(_09992_ ), .B2(_09984_ ), .ZN(_10000_ ) );
AOI21_X1 _13616_ ( .A(fanout_net_11 ), .B1(_09999_ ), .B2(_10000_ ), .ZN(_00238_ ) );
BUF_X4 _13617_ ( .A(_09990_ ), .Z(_10001_ ) );
NAND4_X1 _13618_ ( .A1(_09954_ ), .A2(_09740_ ), .A3(_09931_ ), .A4(_10001_ ), .ZN(_10002_ ) );
OAI21_X1 _13619_ ( .A(\u_lsu.pmem[36] ), .B1(_09992_ ), .B2(_09984_ ), .ZN(_10003_ ) );
AOI21_X1 _13620_ ( .A(fanout_net_11 ), .B1(_10002_ ), .B2(_10003_ ), .ZN(_00239_ ) );
BUF_X4 _13621_ ( .A(_09456_ ), .Z(_10004_ ) );
NAND4_X1 _13622_ ( .A1(_09954_ ), .A2(_10004_ ), .A3(_09934_ ), .A4(_10001_ ), .ZN(_10005_ ) );
OAI21_X1 _13623_ ( .A(\u_lsu.pmem[35] ), .B1(_09992_ ), .B2(_09984_ ), .ZN(_10006_ ) );
AOI21_X1 _13624_ ( .A(fanout_net_11 ), .B1(_10005_ ), .B2(_10006_ ), .ZN(_00240_ ) );
NOR2_X1 _13625_ ( .A1(_09054_ ), .A2(_09557_ ), .ZN(_10007_ ) );
AND2_X1 _13626_ ( .A1(_10007_ ), .A2(_09046_ ), .ZN(_10008_ ) );
BUF_X4 _13627_ ( .A(_08993_ ), .Z(_10009_ ) );
AND2_X2 _13628_ ( .A1(_10008_ ), .A2(_10009_ ), .ZN(_10010_ ) );
AND2_X1 _13629_ ( .A1(_10010_ ), .A2(_09018_ ), .ZN(_10011_ ) );
CLKBUF_X2 _13630_ ( .A(_09493_ ), .Z(_10012_ ) );
AND2_X1 _13631_ ( .A1(_10011_ ), .A2(_10012_ ), .ZN(_10013_ ) );
OAI21_X1 _13632_ ( .A(_09110_ ), .B1(_10013_ ), .B2(\u_lsu.pmem[3943] ), .ZN(_10014_ ) );
AOI21_X1 _13633_ ( .A(_10014_ ), .B1(_09638_ ), .B2(_10013_ ), .ZN(_00241_ ) );
BUF_X4 _13634_ ( .A(_09610_ ), .Z(_10015_ ) );
NAND4_X1 _13635_ ( .A1(_09954_ ), .A2(_10004_ ), .A3(_10015_ ), .A4(_10001_ ), .ZN(_10016_ ) );
OAI21_X1 _13636_ ( .A(\u_lsu.pmem[34] ), .B1(_09992_ ), .B2(_09984_ ), .ZN(_10017_ ) );
AOI21_X1 _13637_ ( .A(fanout_net_11 ), .B1(_10016_ ), .B2(_10017_ ), .ZN(_00242_ ) );
BUF_X4 _13638_ ( .A(_09953_ ), .Z(_10018_ ) );
NAND4_X1 _13639_ ( .A1(_10018_ ), .A2(_10004_ ), .A3(_09941_ ), .A4(_10001_ ), .ZN(_10019_ ) );
OAI21_X1 _13640_ ( .A(\u_lsu.pmem[33] ), .B1(_09992_ ), .B2(_09984_ ), .ZN(_10020_ ) );
AOI21_X1 _13641_ ( .A(fanout_net_11 ), .B1(_10019_ ), .B2(_10020_ ), .ZN(_00243_ ) );
NOR3_X4 _13642_ ( .A1(_09701_ ), .A2(_09785_ ), .A3(_09786_ ), .ZN(_10021_ ) );
NAND4_X1 _13643_ ( .A1(_10021_ ), .A2(_09868_ ), .A3(_09869_ ), .A4(_09998_ ), .ZN(_10022_ ) );
OAI21_X1 _13644_ ( .A(\u_lsu.pmem[32] ), .B1(_09992_ ), .B2(_09984_ ), .ZN(_10023_ ) );
AOI21_X1 _13645_ ( .A(fanout_net_11 ), .B1(_10022_ ), .B2(_10023_ ), .ZN(_00244_ ) );
AOI21_X1 _13646_ ( .A(\u_lsu.pmem[7] ), .B1(_09499_ ), .B2(_09496_ ), .ZN(_10024_ ) );
BUF_X4 _13647_ ( .A(_09955_ ), .Z(_10025_ ) );
AOI211_X1 _13648_ ( .A(fanout_net_11 ), .B(_10024_ ), .C1(_09565_ ), .C2(_10025_ ), .ZN(_00245_ ) );
BUF_X4 _13649_ ( .A(_09108_ ), .Z(_10026_ ) );
OAI21_X1 _13650_ ( .A(_10026_ ), .B1(_10025_ ), .B2(\u_lsu.pmem[6] ), .ZN(_10027_ ) );
AOI21_X1 _13651_ ( .A(_10027_ ), .B1(_09576_ ), .B2(_10025_ ), .ZN(_00246_ ) );
OAI21_X1 _13652_ ( .A(_10026_ ), .B1(_10025_ ), .B2(\u_lsu.pmem[5] ), .ZN(_10028_ ) );
AOI21_X1 _13653_ ( .A(_10028_ ), .B1(_09583_ ), .B2(_10025_ ), .ZN(_00247_ ) );
OAI21_X1 _13654_ ( .A(_10026_ ), .B1(_09955_ ), .B2(\u_lsu.pmem[4] ), .ZN(_10029_ ) );
AOI21_X1 _13655_ ( .A(_10029_ ), .B1(_09146_ ), .B2(_10025_ ), .ZN(_00248_ ) );
OAI21_X1 _13656_ ( .A(_10026_ ), .B1(_09955_ ), .B2(\u_lsu.pmem[3] ), .ZN(_10030_ ) );
AOI21_X1 _13657_ ( .A(_10030_ ), .B1(_09969_ ), .B2(_10025_ ), .ZN(_00249_ ) );
OAI21_X1 _13658_ ( .A(_10026_ ), .B1(_09955_ ), .B2(\u_lsu.pmem[2] ), .ZN(_10031_ ) );
AOI21_X1 _13659_ ( .A(_10031_ ), .B1(_09973_ ), .B2(_10025_ ), .ZN(_00250_ ) );
OAI21_X1 _13660_ ( .A(_10026_ ), .B1(_09955_ ), .B2(\u_lsu.pmem[1] ), .ZN(_10032_ ) );
AOI21_X1 _13661_ ( .A(_10032_ ), .B1(_09977_ ), .B2(_10025_ ), .ZN(_00251_ ) );
BUF_X4 _13662_ ( .A(_09140_ ), .Z(_10033_ ) );
BUF_X4 _13663_ ( .A(_10033_ ), .Z(_10034_ ) );
NAND4_X1 _13664_ ( .A1(_09733_ ), .A2(_09868_ ), .A3(_09869_ ), .A4(_10034_ ), .ZN(_10035_ ) );
BUF_X8 _13665_ ( .A(_09458_ ), .Z(_10036_ ) );
BUF_X4 _13666_ ( .A(_10036_ ), .Z(_10037_ ) );
OAI21_X1 _13667_ ( .A(\u_lsu.pmem[4353] ), .B1(_10037_ ), .B2(_09469_ ), .ZN(_10038_ ) );
AOI21_X1 _13668_ ( .A(fanout_net_11 ), .B1(_10035_ ), .B2(_10038_ ), .ZN(_00252_ ) );
INV_X1 _13669_ ( .A(_10011_ ), .ZN(_10039_ ) );
BUF_X2 _13670_ ( .A(_10039_ ), .Z(_10040_ ) );
BUF_X4 _13671_ ( .A(_09035_ ), .Z(_10041_ ) );
CLKBUF_X2 _13672_ ( .A(_09137_ ), .Z(_10042_ ) );
OR4_X1 _13673_ ( .A1(_09576_ ), .A2(_10040_ ), .A3(_10041_ ), .A4(_10042_ ), .ZN(_10043_ ) );
BUF_X4 _13674_ ( .A(_10040_ ), .Z(_10044_ ) );
CLKBUF_X3 _13675_ ( .A(_09035_ ), .Z(_10045_ ) );
BUF_X4 _13676_ ( .A(_10045_ ), .Z(_10046_ ) );
BUF_X4 _13677_ ( .A(_10046_ ), .Z(_10047_ ) );
OAI21_X1 _13678_ ( .A(\u_lsu.pmem[3942] ), .B1(_10044_ ), .B2(_10047_ ), .ZN(_10048_ ) );
AOI21_X1 _13679_ ( .A(fanout_net_11 ), .B1(_10043_ ), .B2(_10048_ ), .ZN(_00253_ ) );
OAI21_X1 _13680_ ( .A(_10026_ ), .B1(_09955_ ), .B2(\u_lsu.pmem[0] ), .ZN(_10049_ ) );
AOI21_X1 _13681_ ( .A(_10049_ ), .B1(_09497_ ), .B2(_10025_ ), .ZN(_00254_ ) );
BUF_X4 _13682_ ( .A(_09055_ ), .Z(_10050_ ) );
INV_X1 _13683_ ( .A(_09747_ ), .ZN(_10051_ ) );
NOR2_X2 _13684_ ( .A1(_10050_ ), .A2(_10051_ ), .ZN(_10052_ ) );
BUF_X2 _13685_ ( .A(_09046_ ), .Z(_10053_ ) );
AND2_X1 _13686_ ( .A1(_10052_ ), .A2(_10053_ ), .ZN(_10054_ ) );
BUF_X2 _13687_ ( .A(_10009_ ), .Z(_10055_ ) );
AND2_X1 _13688_ ( .A1(_10054_ ), .A2(_10055_ ), .ZN(_10056_ ) );
AND2_X1 _13689_ ( .A1(_10056_ ), .A2(_09491_ ), .ZN(_10057_ ) );
AND2_X1 _13690_ ( .A1(_10057_ ), .A2(_10041_ ), .ZN(_10058_ ) );
OAI21_X1 _13691_ ( .A(_10026_ ), .B1(_10058_ ), .B2(\u_lsu.pmem[8167] ), .ZN(_10059_ ) );
AOI21_X1 _13692_ ( .A(_10059_ ), .B1(_09638_ ), .B2(_10058_ ), .ZN(_00255_ ) );
NAND3_X1 _13693_ ( .A1(_09577_ ), .A2(_09669_ ), .A3(_09754_ ), .ZN(_10060_ ) );
BUF_X4 _13694_ ( .A(_09873_ ), .Z(_10061_ ) );
NOR2_X1 _13695_ ( .A1(_10060_ ), .A2(_10061_ ), .ZN(_10062_ ) );
BUF_X8 _13696_ ( .A(_09875_ ), .Z(_10063_ ) );
BUF_X4 _13697_ ( .A(_10063_ ), .Z(_10064_ ) );
BUF_X4 _13698_ ( .A(_09877_ ), .Z(_10065_ ) );
BUF_X4 _13699_ ( .A(_10065_ ), .Z(_10066_ ) );
NAND4_X1 _13700_ ( .A1(_10062_ ), .A2(_10064_ ), .A3(_10066_ ), .A4(_10034_ ), .ZN(_10067_ ) );
INV_X1 _13701_ ( .A(_10057_ ), .ZN(_10068_ ) );
BUF_X4 _13702_ ( .A(_10068_ ), .Z(_10069_ ) );
BUF_X8 _13703_ ( .A(_09493_ ), .Z(_10070_ ) );
BUF_X4 _13704_ ( .A(_10070_ ), .Z(_10071_ ) );
OAI21_X1 _13705_ ( .A(\u_lsu.pmem[8166] ), .B1(_10069_ ), .B2(_10071_ ), .ZN(_10072_ ) );
AOI21_X1 _13706_ ( .A(fanout_net_11 ), .B1(_10067_ ), .B2(_10072_ ), .ZN(_00256_ ) );
AND3_X1 _13707_ ( .A1(_09584_ ), .A2(_09786_ ), .A3(_09754_ ), .ZN(_10073_ ) );
BUF_X4 _13708_ ( .A(_09536_ ), .Z(_10074_ ) );
AND2_X2 _13709_ ( .A1(_10073_ ), .A2(_10074_ ), .ZN(_10075_ ) );
NAND4_X1 _13710_ ( .A1(_10075_ ), .A2(_10064_ ), .A3(_10066_ ), .A4(_10034_ ), .ZN(_10076_ ) );
OAI21_X1 _13711_ ( .A(\u_lsu.pmem[8165] ), .B1(_10069_ ), .B2(_10071_ ), .ZN(_10077_ ) );
AOI21_X1 _13712_ ( .A(fanout_net_11 ), .B1(_10076_ ), .B2(_10077_ ), .ZN(_00257_ ) );
AND3_X1 _13713_ ( .A1(_09147_ ), .A2(_09786_ ), .A3(_09754_ ), .ZN(_10078_ ) );
AND2_X4 _13714_ ( .A1(_10078_ ), .A2(_10074_ ), .ZN(_10079_ ) );
NAND4_X1 _13715_ ( .A1(_10079_ ), .A2(_10064_ ), .A3(_10066_ ), .A4(_10034_ ), .ZN(_10080_ ) );
BUF_X4 _13716_ ( .A(_10070_ ), .Z(_10081_ ) );
OAI21_X1 _13717_ ( .A(\u_lsu.pmem[8164] ), .B1(_10069_ ), .B2(_10081_ ), .ZN(_10082_ ) );
AOI21_X1 _13718_ ( .A(fanout_net_11 ), .B1(_10080_ ), .B2(_10082_ ), .ZN(_00258_ ) );
AND3_X1 _13719_ ( .A1(_09447_ ), .A2(_09786_ ), .A3(_09754_ ), .ZN(_10083_ ) );
AND2_X2 _13720_ ( .A1(_10083_ ), .A2(_10074_ ), .ZN(_10084_ ) );
NAND4_X1 _13721_ ( .A1(_10084_ ), .A2(_10064_ ), .A3(_10066_ ), .A4(_10034_ ), .ZN(_10085_ ) );
OAI21_X1 _13722_ ( .A(\u_lsu.pmem[8163] ), .B1(_10069_ ), .B2(_10081_ ), .ZN(_10086_ ) );
AOI21_X1 _13723_ ( .A(fanout_net_11 ), .B1(_10085_ ), .B2(_10086_ ), .ZN(_00259_ ) );
AND3_X1 _13724_ ( .A1(_09610_ ), .A2(_09786_ ), .A3(_09747_ ), .ZN(_10087_ ) );
AND2_X2 _13725_ ( .A1(_10087_ ), .A2(_10074_ ), .ZN(_10088_ ) );
BUF_X4 _13726_ ( .A(_10065_ ), .Z(_10089_ ) );
BUF_X4 _13727_ ( .A(_10033_ ), .Z(_10090_ ) );
NAND4_X1 _13728_ ( .A1(_10088_ ), .A2(_10064_ ), .A3(_10089_ ), .A4(_10090_ ), .ZN(_10091_ ) );
OAI21_X1 _13729_ ( .A(\u_lsu.pmem[8162] ), .B1(_10069_ ), .B2(_10081_ ), .ZN(_10092_ ) );
AOI21_X1 _13730_ ( .A(fanout_net_11 ), .B1(_10091_ ), .B2(_10092_ ), .ZN(_00260_ ) );
BUF_X4 _13731_ ( .A(_09873_ ), .Z(_10093_ ) );
NOR3_X4 _13732_ ( .A1(_09783_ ), .A2(_09702_ ), .A3(_10093_ ), .ZN(_10094_ ) );
NAND4_X1 _13733_ ( .A1(_10094_ ), .A2(_10064_ ), .A3(_10089_ ), .A4(_10090_ ), .ZN(_10095_ ) );
OAI21_X1 _13734_ ( .A(\u_lsu.pmem[8161] ), .B1(_10069_ ), .B2(_10081_ ), .ZN(_10096_ ) );
AOI21_X1 _13735_ ( .A(fanout_net_11 ), .B1(_10095_ ), .B2(_10096_ ), .ZN(_00261_ ) );
AND3_X1 _13736_ ( .A1(_09620_ ), .A2(_09786_ ), .A3(_09747_ ), .ZN(_10097_ ) );
AND2_X2 _13737_ ( .A1(_10097_ ), .A2(_10074_ ), .ZN(_10098_ ) );
NAND4_X1 _13738_ ( .A1(_10098_ ), .A2(_10064_ ), .A3(_10089_ ), .A4(_10090_ ), .ZN(_10099_ ) );
OAI21_X1 _13739_ ( .A(\u_lsu.pmem[8160] ), .B1(_10069_ ), .B2(_10081_ ), .ZN(_10100_ ) );
AOI21_X1 _13740_ ( .A(fanout_net_11 ), .B1(_10099_ ), .B2(_10100_ ), .ZN(_00262_ ) );
INV_X1 _13741_ ( .A(_09796_ ), .ZN(_10101_ ) );
NOR2_X2 _13742_ ( .A1(_09463_ ), .A2(_10101_ ), .ZN(_10102_ ) );
AND2_X1 _13743_ ( .A1(_10102_ ), .A2(_09594_ ), .ZN(_10103_ ) );
AND2_X1 _13744_ ( .A1(_10103_ ), .A2(_09489_ ), .ZN(_10104_ ) );
AND2_X1 _13745_ ( .A1(_10104_ ), .A2(_09491_ ), .ZN(_10105_ ) );
INV_X1 _13746_ ( .A(_10105_ ), .ZN(_10106_ ) );
BUF_X4 _13747_ ( .A(_10106_ ), .Z(_10107_ ) );
BUF_X4 _13748_ ( .A(_09496_ ), .Z(_10108_ ) );
OAI21_X1 _13749_ ( .A(\u_lsu.pmem[8135] ), .B1(_10107_ ), .B2(_10108_ ), .ZN(_10109_ ) );
BUF_X4 _13750_ ( .A(_10041_ ), .Z(_10110_ ) );
BUF_X4 _13751_ ( .A(_09605_ ), .Z(_10111_ ) );
NAND4_X1 _13752_ ( .A1(_10104_ ), .A2(_09603_ ), .A3(_10110_ ), .A4(_10111_ ), .ZN(_10112_ ) );
AOI21_X1 _13753_ ( .A(fanout_net_11 ), .B1(_10109_ ), .B2(_10112_ ), .ZN(_00263_ ) );
CLKBUF_X2 _13754_ ( .A(_09035_ ), .Z(_10113_ ) );
OR4_X1 _13755_ ( .A1(_09583_ ), .A2(_10040_ ), .A3(_10113_ ), .A4(_10042_ ), .ZN(_10114_ ) );
OAI21_X1 _13756_ ( .A(\u_lsu.pmem[3941] ), .B1(_10044_ ), .B2(_10047_ ), .ZN(_10115_ ) );
AOI21_X1 _13757_ ( .A(fanout_net_11 ), .B1(_10114_ ), .B2(_10115_ ), .ZN(_00264_ ) );
AND3_X1 _13758_ ( .A1(_09577_ ), .A2(_09668_ ), .A3(_09802_ ), .ZN(_10116_ ) );
AND2_X2 _13759_ ( .A1(_10116_ ), .A2(_10074_ ), .ZN(_10117_ ) );
NAND4_X1 _13760_ ( .A1(_10117_ ), .A2(_10064_ ), .A3(_10089_ ), .A4(_10090_ ), .ZN(_10118_ ) );
OAI21_X1 _13761_ ( .A(\u_lsu.pmem[8134] ), .B1(_10107_ ), .B2(_10081_ ), .ZN(_10119_ ) );
AOI21_X1 _13762_ ( .A(fanout_net_11 ), .B1(_10118_ ), .B2(_10119_ ), .ZN(_00265_ ) );
AND3_X1 _13763_ ( .A1(_09584_ ), .A2(_09668_ ), .A3(_09802_ ), .ZN(_10120_ ) );
AND2_X2 _13764_ ( .A1(_10120_ ), .A2(_10074_ ), .ZN(_10121_ ) );
NAND4_X1 _13765_ ( .A1(_10121_ ), .A2(_10064_ ), .A3(_10089_ ), .A4(_10090_ ), .ZN(_10122_ ) );
OAI21_X1 _13766_ ( .A(\u_lsu.pmem[8133] ), .B1(_10107_ ), .B2(_10081_ ), .ZN(_10123_ ) );
AOI21_X1 _13767_ ( .A(fanout_net_11 ), .B1(_10122_ ), .B2(_10123_ ), .ZN(_00266_ ) );
AND3_X1 _13768_ ( .A1(_09147_ ), .A2(_09668_ ), .A3(_09802_ ), .ZN(_10124_ ) );
AND2_X4 _13769_ ( .A1(_10124_ ), .A2(_10074_ ), .ZN(_10125_ ) );
BUF_X4 _13770_ ( .A(_09875_ ), .Z(_10126_ ) );
BUF_X4 _13771_ ( .A(_10126_ ), .Z(_10127_ ) );
NAND4_X1 _13772_ ( .A1(_10125_ ), .A2(_10127_ ), .A3(_10089_ ), .A4(_10090_ ), .ZN(_10128_ ) );
OAI21_X1 _13773_ ( .A(\u_lsu.pmem[8132] ), .B1(_10107_ ), .B2(_10081_ ), .ZN(_10129_ ) );
AOI21_X1 _13774_ ( .A(fanout_net_11 ), .B1(_10128_ ), .B2(_10129_ ), .ZN(_00267_ ) );
AND3_X1 _13775_ ( .A1(_09447_ ), .A2(_09668_ ), .A3(_09802_ ), .ZN(_10130_ ) );
AND2_X2 _13776_ ( .A1(_10130_ ), .A2(_10074_ ), .ZN(_10131_ ) );
NAND4_X1 _13777_ ( .A1(_10131_ ), .A2(_10127_ ), .A3(_10089_ ), .A4(_10090_ ), .ZN(_10132_ ) );
OAI21_X1 _13778_ ( .A(\u_lsu.pmem[8131] ), .B1(_10107_ ), .B2(_10081_ ), .ZN(_10133_ ) );
AOI21_X1 _13779_ ( .A(fanout_net_11 ), .B1(_10132_ ), .B2(_10133_ ), .ZN(_00268_ ) );
AND3_X1 _13780_ ( .A1(_09610_ ), .A2(_09668_ ), .A3(_09796_ ), .ZN(_10134_ ) );
AND2_X2 _13781_ ( .A1(_10134_ ), .A2(_10074_ ), .ZN(_10135_ ) );
NAND4_X1 _13782_ ( .A1(_10135_ ), .A2(_10127_ ), .A3(_10089_ ), .A4(_10090_ ), .ZN(_10136_ ) );
OAI21_X1 _13783_ ( .A(\u_lsu.pmem[8130] ), .B1(_10107_ ), .B2(_10081_ ), .ZN(_10137_ ) );
AOI21_X1 _13784_ ( .A(fanout_net_11 ), .B1(_10136_ ), .B2(_10137_ ), .ZN(_00269_ ) );
NOR3_X4 _13785_ ( .A1(_09830_ ), .A2(_09702_ ), .A3(_10093_ ), .ZN(_10138_ ) );
NAND4_X1 _13786_ ( .A1(_10138_ ), .A2(_10127_ ), .A3(_10089_ ), .A4(_10090_ ), .ZN(_10139_ ) );
BUF_X4 _13787_ ( .A(_10070_ ), .Z(_10140_ ) );
OAI21_X1 _13788_ ( .A(\u_lsu.pmem[8129] ), .B1(_10107_ ), .B2(_10140_ ), .ZN(_10141_ ) );
AOI21_X1 _13789_ ( .A(fanout_net_11 ), .B1(_10139_ ), .B2(_10141_ ), .ZN(_00270_ ) );
AND3_X1 _13790_ ( .A1(_09620_ ), .A2(_09668_ ), .A3(_09796_ ), .ZN(_10142_ ) );
BUF_X4 _13791_ ( .A(_09536_ ), .Z(_10143_ ) );
AND2_X2 _13792_ ( .A1(_10142_ ), .A2(_10143_ ), .ZN(_10144_ ) );
NAND4_X1 _13793_ ( .A1(_10144_ ), .A2(_10127_ ), .A3(_10089_ ), .A4(_10090_ ), .ZN(_10145_ ) );
OAI21_X1 _13794_ ( .A(\u_lsu.pmem[8128] ), .B1(_10107_ ), .B2(_10140_ ), .ZN(_10146_ ) );
AOI21_X1 _13795_ ( .A(fanout_net_11 ), .B1(_10145_ ), .B2(_10146_ ), .ZN(_00271_ ) );
AND3_X1 _13796_ ( .A1(_09566_ ), .A2(_09668_ ), .A3(_09485_ ), .ZN(_10147_ ) );
AND2_X2 _13797_ ( .A1(_10147_ ), .A2(_10143_ ), .ZN(_10148_ ) );
BUF_X4 _13798_ ( .A(_10065_ ), .Z(_10149_ ) );
BUF_X4 _13799_ ( .A(_10033_ ), .Z(_10150_ ) );
NAND4_X1 _13800_ ( .A1(_10148_ ), .A2(_10127_ ), .A3(_10149_ ), .A4(_10150_ ), .ZN(_10151_ ) );
AND2_X1 _13801_ ( .A1(_09492_ ), .A2(_10045_ ), .ZN(_10152_ ) );
INV_X1 _13802_ ( .A(_10152_ ), .ZN(_10153_ ) );
NAND2_X1 _13803_ ( .A1(_10153_ ), .A2(\u_lsu.pmem[8103] ), .ZN(_10154_ ) );
AOI21_X1 _13804_ ( .A(fanout_net_11 ), .B1(_10151_ ), .B2(_10154_ ), .ZN(_00272_ ) );
NAND3_X1 _13805_ ( .A1(_09577_ ), .A2(_09669_ ), .A3(_09485_ ), .ZN(_10155_ ) );
NOR2_X1 _13806_ ( .A1(_10155_ ), .A2(_10061_ ), .ZN(_10156_ ) );
NAND4_X1 _13807_ ( .A1(_10156_ ), .A2(_10127_ ), .A3(_10149_ ), .A4(_10150_ ), .ZN(_10157_ ) );
NAND2_X1 _13808_ ( .A1(_10153_ ), .A2(\u_lsu.pmem[8102] ), .ZN(_10158_ ) );
AOI21_X1 _13809_ ( .A(fanout_net_12 ), .B1(_10157_ ), .B2(_10158_ ), .ZN(_00273_ ) );
AND3_X1 _13810_ ( .A1(_09584_ ), .A2(_09668_ ), .A3(_09485_ ), .ZN(_10159_ ) );
AND2_X2 _13811_ ( .A1(_10159_ ), .A2(_10143_ ), .ZN(_10160_ ) );
NAND4_X1 _13812_ ( .A1(_10160_ ), .A2(_10127_ ), .A3(_10149_ ), .A4(_10150_ ), .ZN(_10161_ ) );
NAND2_X1 _13813_ ( .A1(_10153_ ), .A2(\u_lsu.pmem[8101] ), .ZN(_10162_ ) );
AOI21_X1 _13814_ ( .A(fanout_net_12 ), .B1(_10161_ ), .B2(_10162_ ), .ZN(_00274_ ) );
OR4_X1 _13815_ ( .A1(_09146_ ), .A2(_10040_ ), .A3(_10113_ ), .A4(_10042_ ), .ZN(_10163_ ) );
OAI21_X1 _13816_ ( .A(\u_lsu.pmem[3940] ), .B1(_10040_ ), .B2(_10047_ ), .ZN(_10164_ ) );
AOI21_X1 _13817_ ( .A(fanout_net_12 ), .B1(_10163_ ), .B2(_10164_ ), .ZN(_00275_ ) );
BUF_X4 _13818_ ( .A(_09486_ ), .Z(_10165_ ) );
AND3_X2 _13819_ ( .A1(_09148_ ), .A2(_10143_ ), .A3(_10165_ ), .ZN(_10166_ ) );
NAND4_X1 _13820_ ( .A1(_10166_ ), .A2(_10127_ ), .A3(_10149_ ), .A4(_10150_ ), .ZN(_10167_ ) );
NAND2_X1 _13821_ ( .A1(_10153_ ), .A2(\u_lsu.pmem[8100] ), .ZN(_10168_ ) );
AOI21_X1 _13822_ ( .A(fanout_net_12 ), .B1(_10167_ ), .B2(_10168_ ), .ZN(_00276_ ) );
AND3_X2 _13823_ ( .A1(_09447_ ), .A2(_10143_ ), .A3(_10165_ ), .ZN(_10169_ ) );
NAND4_X1 _13824_ ( .A1(_10169_ ), .A2(_10127_ ), .A3(_10149_ ), .A4(_10150_ ), .ZN(_10170_ ) );
NAND2_X1 _13825_ ( .A1(_10153_ ), .A2(\u_lsu.pmem[8099] ), .ZN(_10171_ ) );
AOI21_X1 _13826_ ( .A(fanout_net_12 ), .B1(_10170_ ), .B2(_10171_ ), .ZN(_00277_ ) );
AND3_X2 _13827_ ( .A1(_09611_ ), .A2(_10143_ ), .A3(_10165_ ), .ZN(_10172_ ) );
BUF_X4 _13828_ ( .A(_10126_ ), .Z(_10173_ ) );
NAND4_X1 _13829_ ( .A1(_10172_ ), .A2(_10173_ ), .A3(_10149_ ), .A4(_10150_ ), .ZN(_10174_ ) );
NAND2_X1 _13830_ ( .A1(_10153_ ), .A2(\u_lsu.pmem[8098] ), .ZN(_10175_ ) );
AOI21_X1 _13831_ ( .A(fanout_net_12 ), .B1(_10174_ ), .B2(_10175_ ), .ZN(_00278_ ) );
AND3_X2 _13832_ ( .A1(_09615_ ), .A2(_09762_ ), .A3(_10165_ ), .ZN(_10176_ ) );
NAND4_X1 _13833_ ( .A1(_10176_ ), .A2(_10173_ ), .A3(_10149_ ), .A4(_10150_ ), .ZN(_10177_ ) );
NAND2_X1 _13834_ ( .A1(_10153_ ), .A2(\u_lsu.pmem[8097] ), .ZN(_10178_ ) );
AOI21_X1 _13835_ ( .A(fanout_net_12 ), .B1(_10177_ ), .B2(_10178_ ), .ZN(_00279_ ) );
INV_X1 _13836_ ( .A(\u_lsu.pmem[8096] ), .ZN(_10179_ ) );
MUX2_X1 _13837_ ( .A(_10179_ ), .B(_09497_ ), .S(_10152_ ), .Z(_10180_ ) );
NOR2_X1 _13838_ ( .A1(_10180_ ), .A2(fanout_net_12 ), .ZN(_00280_ ) );
OAI21_X1 _13839_ ( .A(\u_lsu.pmem[8071] ), .B1(_09599_ ), .B2(_09444_ ), .ZN(_10181_ ) );
BUF_X4 _13840_ ( .A(_09950_ ), .Z(_10182_ ) );
NAND4_X1 _13841_ ( .A1(_09601_ ), .A2(_09603_ ), .A3(_09659_ ), .A4(_10182_ ), .ZN(_10183_ ) );
AOI21_X1 _13842_ ( .A(fanout_net_12 ), .B1(_10181_ ), .B2(_10183_ ), .ZN(_00281_ ) );
OAI21_X1 _13843_ ( .A(\u_lsu.pmem[8070] ), .B1(_09599_ ), .B2(_09444_ ), .ZN(_10184_ ) );
BUF_X4 _13844_ ( .A(_09575_ ), .Z(_10185_ ) );
NAND4_X1 _13845_ ( .A1(_09601_ ), .A2(_10185_ ), .A3(_09659_ ), .A4(_10182_ ), .ZN(_10186_ ) );
AOI21_X1 _13846_ ( .A(fanout_net_12 ), .B1(_10184_ ), .B2(_10186_ ), .ZN(_00282_ ) );
OAI21_X1 _13847_ ( .A(\u_lsu.pmem[8069] ), .B1(_09598_ ), .B2(_09444_ ), .ZN(_10187_ ) );
BUF_X4 _13848_ ( .A(_09582_ ), .Z(_10188_ ) );
NAND4_X1 _13849_ ( .A1(_09601_ ), .A2(_10188_ ), .A3(_09659_ ), .A4(_10182_ ), .ZN(_10189_ ) );
AOI21_X1 _13850_ ( .A(fanout_net_12 ), .B1(_10187_ ), .B2(_10189_ ), .ZN(_00283_ ) );
BUF_X4 _13851_ ( .A(_09443_ ), .Z(_10190_ ) );
OAI21_X1 _13852_ ( .A(\u_lsu.pmem[8068] ), .B1(_09598_ ), .B2(_10190_ ), .ZN(_10191_ ) );
BUF_X4 _13853_ ( .A(_08605_ ), .Z(_10192_ ) );
NAND4_X1 _13854_ ( .A1(_09601_ ), .A2(_10192_ ), .A3(_09659_ ), .A4(_10182_ ), .ZN(_10193_ ) );
AOI21_X1 _13855_ ( .A(fanout_net_12 ), .B1(_10191_ ), .B2(_10193_ ), .ZN(_00284_ ) );
OAI21_X1 _13856_ ( .A(\u_lsu.pmem[8067] ), .B1(_09598_ ), .B2(_10190_ ), .ZN(_10194_ ) );
NAND4_X1 _13857_ ( .A1(_09601_ ), .A2(_09520_ ), .A3(_10111_ ), .A4(_10182_ ), .ZN(_10195_ ) );
AOI21_X1 _13858_ ( .A(fanout_net_12 ), .B1(_10194_ ), .B2(_10195_ ), .ZN(_00285_ ) );
OR4_X1 _13859_ ( .A1(_09969_ ), .A2(_10040_ ), .A3(_10113_ ), .A4(_10042_ ), .ZN(_10196_ ) );
OAI21_X1 _13860_ ( .A(\u_lsu.pmem[3939] ), .B1(_10040_ ), .B2(_10047_ ), .ZN(_10197_ ) );
AOI21_X1 _13861_ ( .A(fanout_net_12 ), .B1(_10196_ ), .B2(_10197_ ), .ZN(_00286_ ) );
OAI21_X1 _13862_ ( .A(\u_lsu.pmem[8066] ), .B1(_09598_ ), .B2(_10190_ ), .ZN(_10198_ ) );
NAND4_X1 _13863_ ( .A1(_09874_ ), .A2(_09876_ ), .A3(_09879_ ), .A4(_10182_ ), .ZN(_10199_ ) );
AOI21_X1 _13864_ ( .A(fanout_net_12 ), .B1(_10198_ ), .B2(_10199_ ), .ZN(_00287_ ) );
OAI21_X1 _13865_ ( .A(\u_lsu.pmem[8065] ), .B1(_09598_ ), .B2(_10190_ ), .ZN(_10200_ ) );
NAND4_X1 _13866_ ( .A1(_09601_ ), .A2(_09923_ ), .A3(_10111_ ), .A4(_10182_ ), .ZN(_10201_ ) );
AOI21_X1 _13867_ ( .A(fanout_net_12 ), .B1(_10200_ ), .B2(_10201_ ), .ZN(_00288_ ) );
OAI21_X1 _13868_ ( .A(\u_lsu.pmem[8064] ), .B1(_09598_ ), .B2(_10190_ ), .ZN(_10202_ ) );
NAND4_X1 _13869_ ( .A1(_09601_ ), .A2(_09548_ ), .A3(_10111_ ), .A4(_10182_ ), .ZN(_10203_ ) );
AOI21_X1 _13870_ ( .A(fanout_net_12 ), .B1(_10202_ ), .B2(_10203_ ), .ZN(_00289_ ) );
OAI21_X1 _13871_ ( .A(\u_lsu.pmem[8039] ), .B1(_10044_ ), .B2(_10108_ ), .ZN(_10204_ ) );
NAND4_X1 _13872_ ( .A1(_10010_ ), .A2(_09603_ ), .A3(_10110_ ), .A4(_10111_ ), .ZN(_10205_ ) );
AOI21_X1 _13873_ ( .A(fanout_net_12 ), .B1(_10204_ ), .B2(_10205_ ), .ZN(_00290_ ) );
OAI21_X1 _13874_ ( .A(\u_lsu.pmem[8038] ), .B1(_10044_ ), .B2(_10108_ ), .ZN(_10206_ ) );
NAND4_X1 _13875_ ( .A1(_10010_ ), .A2(_10185_ ), .A3(_10110_ ), .A4(_10111_ ), .ZN(_10207_ ) );
AOI21_X1 _13876_ ( .A(fanout_net_12 ), .B1(_10206_ ), .B2(_10207_ ), .ZN(_00291_ ) );
BUF_X4 _13877_ ( .A(_10070_ ), .Z(_10208_ ) );
OAI21_X1 _13878_ ( .A(\u_lsu.pmem[8037] ), .B1(_10044_ ), .B2(_10208_ ), .ZN(_10209_ ) );
NAND4_X1 _13879_ ( .A1(_10010_ ), .A2(_10188_ ), .A3(_10110_ ), .A4(_10111_ ), .ZN(_10210_ ) );
AOI21_X1 _13880_ ( .A(fanout_net_12 ), .B1(_10209_ ), .B2(_10210_ ), .ZN(_00292_ ) );
OAI21_X1 _13881_ ( .A(\u_lsu.pmem[8036] ), .B1(_10044_ ), .B2(_10208_ ), .ZN(_10211_ ) );
BUF_X4 _13882_ ( .A(_10041_ ), .Z(_10212_ ) );
NAND4_X1 _13883_ ( .A1(_10010_ ), .A2(_10192_ ), .A3(_10212_ ), .A4(_10111_ ), .ZN(_10213_ ) );
AOI21_X1 _13884_ ( .A(fanout_net_12 ), .B1(_10211_ ), .B2(_10213_ ), .ZN(_00293_ ) );
OAI21_X1 _13885_ ( .A(\u_lsu.pmem[8035] ), .B1(_10044_ ), .B2(_10208_ ), .ZN(_10214_ ) );
NAND4_X1 _13886_ ( .A1(_10010_ ), .A2(_09520_ ), .A3(_10212_ ), .A4(_10111_ ), .ZN(_10215_ ) );
AOI21_X1 _13887_ ( .A(fanout_net_12 ), .B1(_10214_ ), .B2(_10215_ ), .ZN(_00294_ ) );
OAI21_X1 _13888_ ( .A(\u_lsu.pmem[8034] ), .B1(_10044_ ), .B2(_10208_ ), .ZN(_10216_ ) );
NAND4_X1 _13889_ ( .A1(_10010_ ), .A2(_09474_ ), .A3(_10212_ ), .A4(_10111_ ), .ZN(_10217_ ) );
AOI21_X1 _13890_ ( .A(fanout_net_12 ), .B1(_10216_ ), .B2(_10217_ ), .ZN(_00295_ ) );
OAI21_X1 _13891_ ( .A(\u_lsu.pmem[8033] ), .B1(_10044_ ), .B2(_10208_ ), .ZN(_10218_ ) );
BUF_X4 _13892_ ( .A(_09606_ ), .Z(_10219_ ) );
NAND4_X1 _13893_ ( .A1(_10010_ ), .A2(_09923_ ), .A3(_10212_ ), .A4(_10219_ ), .ZN(_10220_ ) );
AOI21_X1 _13894_ ( .A(fanout_net_12 ), .B1(_10218_ ), .B2(_10220_ ), .ZN(_00296_ ) );
OR4_X1 _13895_ ( .A1(_09973_ ), .A2(_10039_ ), .A3(_10113_ ), .A4(_10042_ ), .ZN(_10221_ ) );
OAI21_X1 _13896_ ( .A(\u_lsu.pmem[3938] ), .B1(_10040_ ), .B2(_10047_ ), .ZN(_10222_ ) );
AOI21_X1 _13897_ ( .A(fanout_net_12 ), .B1(_10221_ ), .B2(_10222_ ), .ZN(_00297_ ) );
OAI21_X1 _13898_ ( .A(\u_lsu.pmem[8032] ), .B1(_10044_ ), .B2(_10208_ ), .ZN(_10223_ ) );
NAND4_X1 _13899_ ( .A1(_10010_ ), .A2(_09548_ ), .A3(_10212_ ), .A4(_10219_ ), .ZN(_10224_ ) );
AOI21_X1 _13900_ ( .A(fanout_net_12 ), .B1(_10223_ ), .B2(_10224_ ), .ZN(_00298_ ) );
NOR2_X1 _13901_ ( .A1(_09054_ ), .A2(_09630_ ), .ZN(_10225_ ) );
AND2_X1 _13902_ ( .A1(_10225_ ), .A2(_09046_ ), .ZN(_10226_ ) );
AND2_X2 _13903_ ( .A1(_10226_ ), .A2(_10009_ ), .ZN(_10227_ ) );
AND2_X1 _13904_ ( .A1(_10227_ ), .A2(_09018_ ), .ZN(_10228_ ) );
INV_X1 _13905_ ( .A(_10228_ ), .ZN(_10229_ ) );
BUF_X2 _13906_ ( .A(_10229_ ), .Z(_10230_ ) );
BUF_X4 _13907_ ( .A(_10230_ ), .Z(_10231_ ) );
OAI21_X1 _13908_ ( .A(\u_lsu.pmem[8007] ), .B1(_10231_ ), .B2(_10208_ ), .ZN(_10232_ ) );
NAND4_X1 _13909_ ( .A1(_10227_ ), .A2(_09603_ ), .A3(_10212_ ), .A4(_10219_ ), .ZN(_10233_ ) );
AOI21_X1 _13910_ ( .A(fanout_net_12 ), .B1(_10232_ ), .B2(_10233_ ), .ZN(_00299_ ) );
OAI21_X1 _13911_ ( .A(\u_lsu.pmem[8006] ), .B1(_10231_ ), .B2(_10208_ ), .ZN(_10234_ ) );
NAND4_X1 _13912_ ( .A1(_10227_ ), .A2(_10185_ ), .A3(_10212_ ), .A4(_10219_ ), .ZN(_10235_ ) );
AOI21_X1 _13913_ ( .A(fanout_net_12 ), .B1(_10234_ ), .B2(_10235_ ), .ZN(_00300_ ) );
OAI21_X1 _13914_ ( .A(\u_lsu.pmem[8005] ), .B1(_10231_ ), .B2(_10208_ ), .ZN(_10236_ ) );
NAND4_X1 _13915_ ( .A1(_10227_ ), .A2(_10188_ ), .A3(_10212_ ), .A4(_10219_ ), .ZN(_10237_ ) );
AOI21_X1 _13916_ ( .A(fanout_net_12 ), .B1(_10236_ ), .B2(_10237_ ), .ZN(_00301_ ) );
OAI21_X1 _13917_ ( .A(\u_lsu.pmem[8004] ), .B1(_10231_ ), .B2(_10208_ ), .ZN(_10238_ ) );
NAND4_X1 _13918_ ( .A1(_10227_ ), .A2(_10192_ ), .A3(_10212_ ), .A4(_10219_ ), .ZN(_10239_ ) );
AOI21_X1 _13919_ ( .A(fanout_net_12 ), .B1(_10238_ ), .B2(_10239_ ), .ZN(_00302_ ) );
BUF_X4 _13920_ ( .A(_10070_ ), .Z(_10240_ ) );
OAI21_X1 _13921_ ( .A(\u_lsu.pmem[8003] ), .B1(_10231_ ), .B2(_10240_ ), .ZN(_10241_ ) );
NAND4_X1 _13922_ ( .A1(_10227_ ), .A2(_09520_ ), .A3(_10212_ ), .A4(_10219_ ), .ZN(_10242_ ) );
AOI21_X1 _13923_ ( .A(fanout_net_13 ), .B1(_10241_ ), .B2(_10242_ ), .ZN(_00303_ ) );
OAI21_X1 _13924_ ( .A(\u_lsu.pmem[8002] ), .B1(_10231_ ), .B2(_10240_ ), .ZN(_10243_ ) );
BUF_X4 _13925_ ( .A(_10041_ ), .Z(_10244_ ) );
NAND4_X1 _13926_ ( .A1(_10227_ ), .A2(_09474_ ), .A3(_10244_ ), .A4(_10219_ ), .ZN(_10245_ ) );
AOI21_X1 _13927_ ( .A(fanout_net_13 ), .B1(_10243_ ), .B2(_10245_ ), .ZN(_00304_ ) );
OAI21_X1 _13928_ ( .A(\u_lsu.pmem[8001] ), .B1(_10231_ ), .B2(_10240_ ), .ZN(_10246_ ) );
NAND4_X1 _13929_ ( .A1(_10227_ ), .A2(_09923_ ), .A3(_10244_ ), .A4(_10219_ ), .ZN(_10247_ ) );
AOI21_X1 _13930_ ( .A(fanout_net_13 ), .B1(_10246_ ), .B2(_10247_ ), .ZN(_00305_ ) );
OAI21_X1 _13931_ ( .A(\u_lsu.pmem[8000] ), .B1(_10231_ ), .B2(_10240_ ), .ZN(_10248_ ) );
NAND4_X1 _13932_ ( .A1(_10227_ ), .A2(_09548_ ), .A3(_10244_ ), .A4(_10219_ ), .ZN(_10249_ ) );
AOI21_X1 _13933_ ( .A(fanout_net_13 ), .B1(_10248_ ), .B2(_10249_ ), .ZN(_00306_ ) );
AND3_X2 _13934_ ( .A1(_09663_ ), .A2(_09669_ ), .A3(_09762_ ), .ZN(_10250_ ) );
NAND4_X1 _13935_ ( .A1(_10250_ ), .A2(_10173_ ), .A3(_10149_ ), .A4(_10150_ ), .ZN(_10251_ ) );
BUF_X2 _13936_ ( .A(_09045_ ), .Z(_10252_ ) );
AND2_X1 _13937_ ( .A1(_09127_ ), .A2(_10252_ ), .ZN(_10253_ ) );
AND2_X1 _13938_ ( .A1(_10253_ ), .A2(_10009_ ), .ZN(_10254_ ) );
AND2_X1 _13939_ ( .A1(_10254_ ), .A2(_09491_ ), .ZN(_10255_ ) );
INV_X1 _13940_ ( .A(_10255_ ), .ZN(_10256_ ) );
BUF_X4 _13941_ ( .A(_10256_ ), .Z(_10257_ ) );
OAI21_X1 _13942_ ( .A(\u_lsu.pmem[7975] ), .B1(_10257_ ), .B2(_10140_ ), .ZN(_10258_ ) );
AOI21_X1 _13943_ ( .A(fanout_net_13 ), .B1(_10251_ ), .B2(_10258_ ), .ZN(_00307_ ) );
OR4_X1 _13944_ ( .A1(_09977_ ), .A2(_10039_ ), .A3(_10113_ ), .A4(_10042_ ), .ZN(_10259_ ) );
OAI21_X1 _13945_ ( .A(\u_lsu.pmem[3937] ), .B1(_10040_ ), .B2(_10047_ ), .ZN(_10260_ ) );
AOI21_X1 _13946_ ( .A(fanout_net_13 ), .B1(_10259_ ), .B2(_10260_ ), .ZN(_00308_ ) );
BUF_X4 _13947_ ( .A(_09481_ ), .Z(_10261_ ) );
BUF_X2 _13948_ ( .A(_10261_ ), .Z(\alu_result_out[5] ) );
NAND2_X1 _13949_ ( .A1(_09680_ ), .A2(\alu_result_out[5] ), .ZN(_10262_ ) );
NOR2_X4 _13950_ ( .A1(_10262_ ), .A2(_10061_ ), .ZN(_10263_ ) );
NAND4_X1 _13951_ ( .A1(_10263_ ), .A2(_10173_ ), .A3(_10149_ ), .A4(_10150_ ), .ZN(_10264_ ) );
OAI21_X1 _13952_ ( .A(\u_lsu.pmem[7974] ), .B1(_10257_ ), .B2(_10140_ ), .ZN(_10265_ ) );
AOI21_X1 _13953_ ( .A(fanout_net_13 ), .B1(_10264_ ), .B2(_10265_ ), .ZN(_00309_ ) );
NAND2_X1 _13954_ ( .A1(_09684_ ), .A2(\alu_result_out[5] ), .ZN(_10266_ ) );
NOR2_X4 _13955_ ( .A1(_10266_ ), .A2(_10061_ ), .ZN(_10267_ ) );
NAND4_X1 _13956_ ( .A1(_10267_ ), .A2(_10173_ ), .A3(_10149_ ), .A4(_10150_ ), .ZN(_10268_ ) );
OAI21_X1 _13957_ ( .A(\u_lsu.pmem[7973] ), .B1(_10257_ ), .B2(_10140_ ), .ZN(_10269_ ) );
AOI21_X1 _13958_ ( .A(fanout_net_13 ), .B1(_10268_ ), .B2(_10269_ ), .ZN(_00310_ ) );
AND2_X1 _13959_ ( .A1(_09141_ ), .A2(_10255_ ), .ZN(_10270_ ) );
OAI21_X1 _13960_ ( .A(_10026_ ), .B1(_10270_ ), .B2(\u_lsu.pmem[7972] ), .ZN(_10271_ ) );
AOI21_X1 _13961_ ( .A(_10271_ ), .B1(_09691_ ), .B2(_10270_ ), .ZN(_00311_ ) );
OAI21_X1 _13962_ ( .A(\u_lsu.pmem[7971] ), .B1(_10257_ ), .B2(_10240_ ), .ZN(_10272_ ) );
BUF_X4 _13963_ ( .A(_09606_ ), .Z(_10273_ ) );
NAND4_X1 _13964_ ( .A1(_10254_ ), .A2(_09520_ ), .A3(_10244_ ), .A4(_10273_ ), .ZN(_10274_ ) );
AOI21_X1 _13965_ ( .A(fanout_net_13 ), .B1(_10272_ ), .B2(_10274_ ), .ZN(_00312_ ) );
OAI21_X1 _13966_ ( .A(\u_lsu.pmem[7970] ), .B1(_10257_ ), .B2(_10240_ ), .ZN(_10275_ ) );
NAND4_X1 _13967_ ( .A1(_10254_ ), .A2(_09474_ ), .A3(_10244_ ), .A4(_10273_ ), .ZN(_10276_ ) );
AOI21_X1 _13968_ ( .A(fanout_net_13 ), .B1(_10275_ ), .B2(_10276_ ), .ZN(_00313_ ) );
OAI21_X1 _13969_ ( .A(\u_lsu.pmem[7969] ), .B1(_10257_ ), .B2(_10240_ ), .ZN(_10277_ ) );
NAND4_X1 _13970_ ( .A1(_10254_ ), .A2(_09923_ ), .A3(_10244_ ), .A4(_10273_ ), .ZN(_10278_ ) );
AOI21_X1 _13971_ ( .A(fanout_net_13 ), .B1(_10277_ ), .B2(_10278_ ), .ZN(_00314_ ) );
NOR3_X4 _13972_ ( .A1(_09701_ ), .A2(_09535_ ), .A3(_09873_ ), .ZN(_10279_ ) );
BUF_X4 _13973_ ( .A(_10065_ ), .Z(_10280_ ) );
BUF_X4 _13974_ ( .A(_10033_ ), .Z(_10281_ ) );
NAND4_X1 _13975_ ( .A1(_10279_ ), .A2(_10173_ ), .A3(_10280_ ), .A4(_10281_ ), .ZN(_10282_ ) );
OAI21_X1 _13976_ ( .A(\u_lsu.pmem[7968] ), .B1(_10257_ ), .B2(_10140_ ), .ZN(_10283_ ) );
AOI21_X1 _13977_ ( .A(fanout_net_13 ), .B1(_10282_ ), .B2(_10283_ ), .ZN(_00315_ ) );
AND2_X1 _13978_ ( .A1(_09566_ ), .A2(_09707_ ), .ZN(_10284_ ) );
AND2_X2 _13979_ ( .A1(_10284_ ), .A2(\alu_result_out[6] ), .ZN(_10285_ ) );
BUF_X4 _13980_ ( .A(_09489_ ), .Z(_10286_ ) );
BUF_X8 _13981_ ( .A(_10286_ ), .Z(_10287_ ) );
BUF_X2 _13982_ ( .A(_10287_ ), .Z(\alu_result_out[7] ) );
NAND4_X1 _13983_ ( .A1(_10285_ ), .A2(\alu_result_out[7] ), .A3(_10280_ ), .A4(_10281_ ), .ZN(_10288_ ) );
AND2_X1 _13984_ ( .A1(_09465_ ), .A2(_09784_ ), .ZN(_10289_ ) );
AND2_X1 _13985_ ( .A1(_10289_ ), .A2(_10286_ ), .ZN(_10290_ ) );
AND2_X1 _13986_ ( .A1(_10290_ ), .A2(_09605_ ), .ZN(_10291_ ) );
NAND2_X1 _13987_ ( .A1(_09950_ ), .A2(_10291_ ), .ZN(_10292_ ) );
NAND2_X1 _13988_ ( .A1(_10292_ ), .A2(\u_lsu.pmem[7943] ), .ZN(_10293_ ) );
AOI21_X1 _13989_ ( .A(fanout_net_13 ), .B1(_10288_ ), .B2(_10293_ ), .ZN(_00316_ ) );
AND2_X1 _13990_ ( .A1(_09578_ ), .A2(_09707_ ), .ZN(_10294_ ) );
AND2_X2 _13991_ ( .A1(_10294_ ), .A2(\alu_result_out[6] ), .ZN(_10295_ ) );
NAND4_X1 _13992_ ( .A1(_10295_ ), .A2(\alu_result_out[7] ), .A3(_10280_ ), .A4(_10281_ ), .ZN(_10296_ ) );
NAND2_X1 _13993_ ( .A1(_10292_ ), .A2(\u_lsu.pmem[7942] ), .ZN(_10297_ ) );
AOI21_X1 _13994_ ( .A(fanout_net_13 ), .B1(_10296_ ), .B2(_10297_ ), .ZN(_00317_ ) );
AND2_X1 _13995_ ( .A1(_09585_ ), .A2(_09707_ ), .ZN(_10298_ ) );
AND2_X2 _13996_ ( .A1(_10298_ ), .A2(\alu_result_out[6] ), .ZN(_10299_ ) );
NAND4_X1 _13997_ ( .A1(_10299_ ), .A2(\alu_result_out[7] ), .A3(_10280_ ), .A4(_10281_ ), .ZN(_10300_ ) );
NAND2_X1 _13998_ ( .A1(_10292_ ), .A2(\u_lsu.pmem[7941] ), .ZN(_10301_ ) );
AOI21_X1 _13999_ ( .A(fanout_net_13 ), .B1(_10300_ ), .B2(_10301_ ), .ZN(_00318_ ) );
CLKBUF_X2 _14000_ ( .A(_09137_ ), .Z(_10302_ ) );
OR4_X1 _14001_ ( .A1(_09497_ ), .A2(_10039_ ), .A3(_10113_ ), .A4(_10302_ ), .ZN(_10303_ ) );
OAI21_X1 _14002_ ( .A(\u_lsu.pmem[3936] ), .B1(_10040_ ), .B2(_10047_ ), .ZN(_10304_ ) );
AOI21_X1 _14003_ ( .A(fanout_net_13 ), .B1(_10303_ ), .B2(_10304_ ), .ZN(_00319_ ) );
AND2_X1 _14004_ ( .A1(_09147_ ), .A2(_09707_ ), .ZN(_10305_ ) );
AND2_X2 _14005_ ( .A1(_10305_ ), .A2(\alu_result_out[6] ), .ZN(_10306_ ) );
NAND4_X1 _14006_ ( .A1(_10306_ ), .A2(\alu_result_out[7] ), .A3(_10280_ ), .A4(_10281_ ), .ZN(_10307_ ) );
NAND2_X1 _14007_ ( .A1(_10292_ ), .A2(\u_lsu.pmem[7940] ), .ZN(_10308_ ) );
AOI21_X1 _14008_ ( .A(fanout_net_13 ), .B1(_10307_ ), .B2(_10308_ ), .ZN(_00320_ ) );
AND2_X2 _14009_ ( .A1(_09724_ ), .A2(\alu_result_out[6] ), .ZN(_10309_ ) );
NAND4_X1 _14010_ ( .A1(_10309_ ), .A2(\alu_result_out[7] ), .A3(_10280_ ), .A4(_10281_ ), .ZN(_10310_ ) );
NAND2_X1 _14011_ ( .A1(_10292_ ), .A2(\u_lsu.pmem[7939] ), .ZN(_10311_ ) );
AOI21_X1 _14012_ ( .A(fanout_net_13 ), .B1(_10310_ ), .B2(_10311_ ), .ZN(_00321_ ) );
NAND2_X1 _14013_ ( .A1(_10292_ ), .A2(\u_lsu.pmem[7938] ), .ZN(_10312_ ) );
NOR3_X1 _14014_ ( .A1(_09873_ ), .A2(_08962_ ), .A3(_09466_ ), .ZN(_10313_ ) );
NAND4_X1 _14015_ ( .A1(_09473_ ), .A2(_09876_ ), .A3(_09879_ ), .A4(_10313_ ), .ZN(_10314_ ) );
AOI21_X1 _14016_ ( .A(fanout_net_13 ), .B1(_10312_ ), .B2(_10314_ ), .ZN(_00322_ ) );
AND2_X1 _14017_ ( .A1(_09615_ ), .A2(_09465_ ), .ZN(_10315_ ) );
AND2_X2 _14018_ ( .A1(_10315_ ), .A2(\alu_result_out[6] ), .ZN(_10316_ ) );
NAND4_X1 _14019_ ( .A1(_10316_ ), .A2(\alu_result_out[7] ), .A3(_10280_ ), .A4(_10281_ ), .ZN(_10317_ ) );
NAND2_X1 _14020_ ( .A1(_10292_ ), .A2(\u_lsu.pmem[7937] ), .ZN(_10318_ ) );
AOI21_X1 _14021_ ( .A(fanout_net_13 ), .B1(_10317_ ), .B2(_10318_ ), .ZN(_00323_ ) );
AND2_X1 _14022_ ( .A1(_09620_ ), .A2(_09465_ ), .ZN(_10319_ ) );
AND2_X2 _14023_ ( .A1(_10319_ ), .A2(\alu_result_out[6] ), .ZN(_10320_ ) );
NAND4_X1 _14024_ ( .A1(_10320_ ), .A2(\alu_result_out[7] ), .A3(_10280_ ), .A4(_10281_ ), .ZN(_10321_ ) );
NAND2_X1 _14025_ ( .A1(_10292_ ), .A2(\u_lsu.pmem[7936] ), .ZN(_10322_ ) );
AOI21_X1 _14026_ ( .A(fanout_net_13 ), .B1(_10321_ ), .B2(_10322_ ), .ZN(_00324_ ) );
NAND3_X1 _14027_ ( .A1(_09462_ ), .A2(_09744_ ), .A3(_09747_ ), .ZN(_10323_ ) );
NOR2_X1 _14028_ ( .A1(_09506_ ), .A2(_10323_ ), .ZN(_10324_ ) );
BUF_X4 _14029_ ( .A(_09134_ ), .Z(_10325_ ) );
BUF_X4 _14030_ ( .A(_10325_ ), .Z(_10326_ ) );
NAND2_X1 _14031_ ( .A1(_10324_ ), .A2(_10326_ ), .ZN(_10327_ ) );
BUF_X4 _14032_ ( .A(_10327_ ), .Z(_10328_ ) );
OAI21_X1 _14033_ ( .A(\u_lsu.pmem[7911] ), .B1(_09460_ ), .B2(_10328_ ), .ZN(_10329_ ) );
BUF_X4 _14034_ ( .A(_09741_ ), .Z(_10330_ ) );
NAND4_X1 _14035_ ( .A1(_10330_ ), .A2(_09452_ ), .A3(_09879_ ), .A4(_10324_ ), .ZN(_10331_ ) );
AOI21_X1 _14036_ ( .A(fanout_net_13 ), .B1(_10329_ ), .B2(_10331_ ), .ZN(_00325_ ) );
AND2_X2 _14037_ ( .A1(_09755_ ), .A2(_10143_ ), .ZN(_10332_ ) );
NAND4_X1 _14038_ ( .A1(_10332_ ), .A2(_10173_ ), .A3(_10280_ ), .A4(_10281_ ), .ZN(_10333_ ) );
BUF_X4 _14039_ ( .A(_10036_ ), .Z(_10334_ ) );
OAI21_X1 _14040_ ( .A(\u_lsu.pmem[7910] ), .B1(_10334_ ), .B2(_10328_ ), .ZN(_10335_ ) );
AOI21_X1 _14041_ ( .A(fanout_net_13 ), .B1(_10333_ ), .B2(_10335_ ), .ZN(_00326_ ) );
NOR2_X1 _14042_ ( .A1(_09761_ ), .A2(_10061_ ), .ZN(_10336_ ) );
NAND4_X1 _14043_ ( .A1(_10336_ ), .A2(_10173_ ), .A3(_10280_ ), .A4(_10281_ ), .ZN(_10337_ ) );
OAI21_X1 _14044_ ( .A(\u_lsu.pmem[7909] ), .B1(_10334_ ), .B2(_10328_ ), .ZN(_10338_ ) );
AOI21_X1 _14045_ ( .A(fanout_net_13 ), .B1(_10337_ ), .B2(_10338_ ), .ZN(_00327_ ) );
AND2_X4 _14046_ ( .A1(_09769_ ), .A2(_10143_ ), .ZN(_10339_ ) );
BUF_X8 _14047_ ( .A(_09877_ ), .Z(_10340_ ) );
BUF_X4 _14048_ ( .A(_10340_ ), .Z(_10341_ ) );
BUF_X4 _14049_ ( .A(_10033_ ), .Z(_10342_ ) );
NAND4_X1 _14050_ ( .A1(_10339_ ), .A2(_10173_ ), .A3(_10341_ ), .A4(_10342_ ), .ZN(_10343_ ) );
OAI21_X1 _14051_ ( .A(\u_lsu.pmem[7908] ), .B1(_10334_ ), .B2(_10328_ ), .ZN(_10344_ ) );
AOI21_X1 _14052_ ( .A(fanout_net_13 ), .B1(_10343_ ), .B2(_10344_ ), .ZN(_00328_ ) );
NOR2_X2 _14053_ ( .A1(_09773_ ), .A2(_10061_ ), .ZN(_10345_ ) );
NAND4_X1 _14054_ ( .A1(_10345_ ), .A2(_10173_ ), .A3(_10341_ ), .A4(_10342_ ), .ZN(_10346_ ) );
OAI21_X1 _14055_ ( .A(\u_lsu.pmem[7907] ), .B1(_10334_ ), .B2(_10328_ ), .ZN(_10347_ ) );
AOI21_X1 _14056_ ( .A(fanout_net_13 ), .B1(_10346_ ), .B2(_10347_ ), .ZN(_00329_ ) );
AND2_X1 _14057_ ( .A1(_10228_ ), .A2(_10012_ ), .ZN(_10348_ ) );
OAI21_X1 _14058_ ( .A(_10026_ ), .B1(_10348_ ), .B2(\u_lsu.pmem[3911] ), .ZN(_10349_ ) );
AOI21_X1 _14059_ ( .A(_10349_ ), .B1(_09638_ ), .B2(_10348_ ), .ZN(_00330_ ) );
NOR2_X4 _14060_ ( .A1(_09779_ ), .A2(_10061_ ), .ZN(_10350_ ) );
BUF_X4 _14061_ ( .A(_10126_ ), .Z(_10351_ ) );
NAND4_X1 _14062_ ( .A1(_10350_ ), .A2(_10351_ ), .A3(_10341_ ), .A4(_10342_ ), .ZN(_10352_ ) );
OAI21_X1 _14063_ ( .A(\u_lsu.pmem[7906] ), .B1(_10334_ ), .B2(_10328_ ), .ZN(_10353_ ) );
AOI21_X1 _14064_ ( .A(fanout_net_13 ), .B1(_10352_ ), .B2(_10353_ ), .ZN(_00331_ ) );
NOR3_X4 _14065_ ( .A1(_09783_ ), .A2(_09669_ ), .A3(_09873_ ), .ZN(_10354_ ) );
NAND4_X1 _14066_ ( .A1(_10354_ ), .A2(_10351_ ), .A3(_10341_ ), .A4(_10342_ ), .ZN(_10355_ ) );
OAI21_X1 _14067_ ( .A(\u_lsu.pmem[7905] ), .B1(_10334_ ), .B2(_10328_ ), .ZN(_10356_ ) );
AOI21_X1 _14068_ ( .A(fanout_net_13 ), .B1(_10355_ ), .B2(_10356_ ), .ZN(_00332_ ) );
NOR2_X2 _14069_ ( .A1(_09790_ ), .A2(_10061_ ), .ZN(_10357_ ) );
NAND4_X1 _14070_ ( .A1(_10357_ ), .A2(_10351_ ), .A3(_10341_ ), .A4(_10342_ ), .ZN(_10358_ ) );
OAI21_X1 _14071_ ( .A(\u_lsu.pmem[7904] ), .B1(_10334_ ), .B2(_10328_ ), .ZN(_10359_ ) );
AOI21_X1 _14072_ ( .A(fanout_net_13 ), .B1(_10358_ ), .B2(_10359_ ), .ZN(_00333_ ) );
BUF_X4 _14073_ ( .A(_09572_ ), .Z(_10360_ ) );
NAND3_X1 _14074_ ( .A1(_09462_ ), .A2(_09744_ ), .A3(_09796_ ), .ZN(_10361_ ) );
NOR2_X1 _14075_ ( .A1(_09506_ ), .A2(_10361_ ), .ZN(_10362_ ) );
NAND2_X1 _14076_ ( .A1(_10362_ ), .A2(_10326_ ), .ZN(_10363_ ) );
BUF_X4 _14077_ ( .A(_10363_ ), .Z(_10364_ ) );
OAI21_X1 _14078_ ( .A(\u_lsu.pmem[7879] ), .B1(_10360_ ), .B2(_10364_ ), .ZN(_10365_ ) );
BUF_X4 _14079_ ( .A(_09451_ ), .Z(_10366_ ) );
NAND4_X1 _14080_ ( .A1(_10330_ ), .A2(_10366_ ), .A3(_09879_ ), .A4(_10362_ ), .ZN(_10367_ ) );
AOI21_X1 _14081_ ( .A(fanout_net_13 ), .B1(_10365_ ), .B2(_10367_ ), .ZN(_00334_ ) );
NOR2_X4 _14082_ ( .A1(_09803_ ), .A2(_10061_ ), .ZN(_10368_ ) );
NAND4_X1 _14083_ ( .A1(_10368_ ), .A2(_10351_ ), .A3(_10341_ ), .A4(_10342_ ), .ZN(_10369_ ) );
OAI21_X1 _14084_ ( .A(\u_lsu.pmem[7878] ), .B1(_10334_ ), .B2(_10364_ ), .ZN(_10370_ ) );
AOI21_X1 _14085_ ( .A(fanout_net_14 ), .B1(_10369_ ), .B2(_10370_ ), .ZN(_00335_ ) );
NOR2_X1 _14086_ ( .A1(_09810_ ), .A2(_10093_ ), .ZN(_10371_ ) );
NAND4_X1 _14087_ ( .A1(_10371_ ), .A2(_10351_ ), .A3(_10341_ ), .A4(_10342_ ), .ZN(_10372_ ) );
OAI21_X1 _14088_ ( .A(\u_lsu.pmem[7877] ), .B1(_10334_ ), .B2(_10364_ ), .ZN(_10373_ ) );
AOI21_X1 _14089_ ( .A(fanout_net_14 ), .B1(_10372_ ), .B2(_10373_ ), .ZN(_00336_ ) );
AND2_X4 _14090_ ( .A1(_09814_ ), .A2(_10143_ ), .ZN(_10374_ ) );
NAND4_X1 _14091_ ( .A1(_10374_ ), .A2(_10351_ ), .A3(_10341_ ), .A4(_10342_ ), .ZN(_10375_ ) );
OAI21_X1 _14092_ ( .A(\u_lsu.pmem[7876] ), .B1(_10334_ ), .B2(_10364_ ), .ZN(_10376_ ) );
AOI21_X1 _14093_ ( .A(fanout_net_14 ), .B1(_10375_ ), .B2(_10376_ ), .ZN(_00337_ ) );
AND2_X2 _14094_ ( .A1(_09818_ ), .A2(_10143_ ), .ZN(_10377_ ) );
NAND4_X1 _14095_ ( .A1(_10377_ ), .A2(_10351_ ), .A3(_10341_ ), .A4(_10342_ ), .ZN(_10378_ ) );
BUF_X4 _14096_ ( .A(_10036_ ), .Z(_10379_ ) );
OAI21_X1 _14097_ ( .A(\u_lsu.pmem[7875] ), .B1(_10379_ ), .B2(_10364_ ), .ZN(_10380_ ) );
AOI21_X1 _14098_ ( .A(fanout_net_14 ), .B1(_10378_ ), .B2(_10380_ ), .ZN(_00338_ ) );
NOR2_X4 _14099_ ( .A1(_09826_ ), .A2(_10093_ ), .ZN(_10381_ ) );
NAND4_X1 _14100_ ( .A1(_10381_ ), .A2(_10351_ ), .A3(_10341_ ), .A4(_10342_ ), .ZN(_10382_ ) );
OAI21_X1 _14101_ ( .A(\u_lsu.pmem[7874] ), .B1(_10379_ ), .B2(_10364_ ), .ZN(_10383_ ) );
AOI21_X1 _14102_ ( .A(fanout_net_14 ), .B1(_10382_ ), .B2(_10383_ ), .ZN(_00339_ ) );
NOR3_X4 _14103_ ( .A1(_09830_ ), .A2(_09669_ ), .A3(_09873_ ), .ZN(_10384_ ) );
BUF_X4 _14104_ ( .A(_10340_ ), .Z(_10385_ ) );
BUF_X4 _14105_ ( .A(_10033_ ), .Z(_10386_ ) );
NAND4_X1 _14106_ ( .A1(_10384_ ), .A2(_10351_ ), .A3(_10385_ ), .A4(_10386_ ), .ZN(_10387_ ) );
OAI21_X1 _14107_ ( .A(\u_lsu.pmem[7873] ), .B1(_10379_ ), .B2(_10364_ ), .ZN(_10388_ ) );
AOI21_X1 _14108_ ( .A(fanout_net_14 ), .B1(_10387_ ), .B2(_10388_ ), .ZN(_00340_ ) );
OR4_X1 _14109_ ( .A1(_09576_ ), .A2(_10230_ ), .A3(_10113_ ), .A4(_10302_ ), .ZN(_10389_ ) );
OAI21_X1 _14110_ ( .A(\u_lsu.pmem[3910] ), .B1(_10231_ ), .B2(_10047_ ), .ZN(_10390_ ) );
AOI21_X1 _14111_ ( .A(fanout_net_14 ), .B1(_10389_ ), .B2(_10390_ ), .ZN(_00341_ ) );
NOR2_X2 _14112_ ( .A1(_09834_ ), .A2(_10093_ ), .ZN(_10391_ ) );
NAND4_X1 _14113_ ( .A1(_10391_ ), .A2(_10351_ ), .A3(_10385_ ), .A4(_10386_ ), .ZN(_10392_ ) );
OAI21_X1 _14114_ ( .A(\u_lsu.pmem[7872] ), .B1(_10379_ ), .B2(_10364_ ), .ZN(_10393_ ) );
AOI21_X1 _14115_ ( .A(fanout_net_14 ), .B1(_10392_ ), .B2(_10393_ ), .ZN(_00342_ ) );
NOR2_X1 _14116_ ( .A1(_09839_ ), .A2(_10093_ ), .ZN(_10394_ ) );
BUF_X4 _14117_ ( .A(_10126_ ), .Z(_10395_ ) );
NAND4_X1 _14118_ ( .A1(_10394_ ), .A2(_10395_ ), .A3(_10385_ ), .A4(_10386_ ), .ZN(_10396_ ) );
BUF_X4 _14119_ ( .A(_09118_ ), .Z(_10397_ ) );
AND3_X2 _14120_ ( .A1(_10397_ ), .A2(_09462_ ), .A3(_09857_ ), .ZN(_10398_ ) );
NAND2_X1 _14121_ ( .A1(_10398_ ), .A2(_10326_ ), .ZN(_10399_ ) );
BUF_X4 _14122_ ( .A(_10399_ ), .Z(_10400_ ) );
OAI21_X1 _14123_ ( .A(\u_lsu.pmem[7847] ), .B1(_10379_ ), .B2(_10400_ ), .ZN(_10401_ ) );
AOI21_X1 _14124_ ( .A(fanout_net_14 ), .B1(_10396_ ), .B2(_10401_ ), .ZN(_00343_ ) );
NOR2_X1 _14125_ ( .A1(_09848_ ), .A2(_10093_ ), .ZN(_10402_ ) );
NAND4_X1 _14126_ ( .A1(_10402_ ), .A2(_10395_ ), .A3(_10385_ ), .A4(_10386_ ), .ZN(_10403_ ) );
OAI21_X1 _14127_ ( .A(\u_lsu.pmem[7846] ), .B1(_10379_ ), .B2(_10400_ ), .ZN(_10404_ ) );
AOI21_X1 _14128_ ( .A(fanout_net_14 ), .B1(_10403_ ), .B2(_10404_ ), .ZN(_00344_ ) );
NOR2_X1 _14129_ ( .A1(_09852_ ), .A2(_10093_ ), .ZN(_10405_ ) );
NAND4_X1 _14130_ ( .A1(_10405_ ), .A2(_10395_ ), .A3(_10385_ ), .A4(_10386_ ), .ZN(_10406_ ) );
OAI21_X1 _14131_ ( .A(\u_lsu.pmem[7845] ), .B1(_10379_ ), .B2(_10400_ ), .ZN(_10407_ ) );
AOI21_X1 _14132_ ( .A(fanout_net_14 ), .B1(_10406_ ), .B2(_10407_ ), .ZN(_00345_ ) );
AND3_X2 _14133_ ( .A1(_09148_ ), .A2(_09762_ ), .A3(_09857_ ), .ZN(_10408_ ) );
NAND4_X1 _14134_ ( .A1(_10408_ ), .A2(_10395_ ), .A3(_10385_ ), .A4(_10386_ ), .ZN(_10409_ ) );
OAI21_X1 _14135_ ( .A(\u_lsu.pmem[7844] ), .B1(_10379_ ), .B2(_10400_ ), .ZN(_10410_ ) );
AOI21_X1 _14136_ ( .A(fanout_net_14 ), .B1(_10409_ ), .B2(_10410_ ), .ZN(_00346_ ) );
AND3_X2 _14137_ ( .A1(_09447_ ), .A2(_09762_ ), .A3(_09857_ ), .ZN(_10411_ ) );
NAND4_X1 _14138_ ( .A1(_10411_ ), .A2(_10395_ ), .A3(_10385_ ), .A4(_10386_ ), .ZN(_10412_ ) );
OAI21_X1 _14139_ ( .A(\u_lsu.pmem[7843] ), .B1(_10379_ ), .B2(_10400_ ), .ZN(_10413_ ) );
AOI21_X1 _14140_ ( .A(fanout_net_14 ), .B1(_10412_ ), .B2(_10413_ ), .ZN(_00347_ ) );
AND3_X2 _14141_ ( .A1(_09611_ ), .A2(_09762_ ), .A3(_09857_ ), .ZN(_10414_ ) );
NAND4_X1 _14142_ ( .A1(_10414_ ), .A2(_10395_ ), .A3(_10385_ ), .A4(_10386_ ), .ZN(_10415_ ) );
OAI21_X1 _14143_ ( .A(\u_lsu.pmem[7842] ), .B1(_10379_ ), .B2(_10400_ ), .ZN(_10416_ ) );
AOI21_X1 _14144_ ( .A(fanout_net_14 ), .B1(_10415_ ), .B2(_10416_ ), .ZN(_00348_ ) );
AND3_X2 _14145_ ( .A1(_09615_ ), .A2(_09762_ ), .A3(_09857_ ), .ZN(_10417_ ) );
NAND4_X1 _14146_ ( .A1(_10417_ ), .A2(_10395_ ), .A3(_10385_ ), .A4(_10386_ ), .ZN(_10418_ ) );
BUF_X4 _14147_ ( .A(_10036_ ), .Z(_10419_ ) );
OAI21_X1 _14148_ ( .A(\u_lsu.pmem[7841] ), .B1(_10419_ ), .B2(_10400_ ), .ZN(_10420_ ) );
AOI21_X1 _14149_ ( .A(fanout_net_14 ), .B1(_10418_ ), .B2(_10420_ ), .ZN(_00349_ ) );
OAI21_X1 _14150_ ( .A(\u_lsu.pmem[7840] ), .B1(_10360_ ), .B2(_10400_ ), .ZN(_10421_ ) );
NAND4_X1 _14151_ ( .A1(_09622_ ), .A2(_10366_ ), .A3(_09879_ ), .A4(_10398_ ), .ZN(_10422_ ) );
AOI21_X1 _14152_ ( .A(fanout_net_14 ), .B1(_10421_ ), .B2(_10422_ ), .ZN(_00350_ ) );
AND3_X2 _14153_ ( .A1(_09503_ ), .A2(_09534_ ), .A3(_09462_ ), .ZN(_10423_ ) );
BUF_X4 _14154_ ( .A(_09134_ ), .Z(_10424_ ) );
NAND3_X1 _14155_ ( .A1(_10423_ ), .A2(_09875_ ), .A3(_10424_ ), .ZN(_10425_ ) );
BUF_X4 _14156_ ( .A(_10425_ ), .Z(_10426_ ) );
OAI21_X1 _14157_ ( .A(\u_lsu.pmem[7815] ), .B1(_10426_ ), .B2(_10190_ ), .ZN(_10427_ ) );
INV_X1 _14158_ ( .A(_09066_ ), .ZN(_10428_ ) );
CLKBUF_X3 _14159_ ( .A(_10428_ ), .Z(_10429_ ) );
BUF_X2 _14160_ ( .A(_10429_ ), .Z(_10430_ ) );
BUF_X4 _14161_ ( .A(_10430_ ), .Z(_10431_ ) );
BUF_X4 _14162_ ( .A(_10431_ ), .Z(_10432_ ) );
BUF_X4 _14163_ ( .A(_10432_ ), .Z(_10433_ ) );
AND3_X1 _14164_ ( .A1(_09566_ ), .A2(_10433_ ), .A3(_09096_ ), .ZN(_10434_ ) );
NAND3_X1 _14165_ ( .A1(_10434_ ), .A2(_09888_ ), .A3(_09532_ ), .ZN(_10435_ ) );
NOR2_X4 _14166_ ( .A1(_10435_ ), .A2(_10093_ ), .ZN(_10436_ ) );
BUF_X4 _14167_ ( .A(_10063_ ), .Z(_10437_ ) );
BUF_X4 _14168_ ( .A(_09878_ ), .Z(_10438_ ) );
NAND4_X1 _14169_ ( .A1(_10436_ ), .A2(_10437_ ), .A3(_10438_ ), .A4(_10182_ ), .ZN(_10439_ ) );
AOI21_X1 _14170_ ( .A(fanout_net_14 ), .B1(_10427_ ), .B2(_10439_ ), .ZN(_00351_ ) );
OR4_X1 _14171_ ( .A1(_09583_ ), .A2(_10230_ ), .A3(_10113_ ), .A4(_10302_ ), .ZN(_10440_ ) );
OAI21_X1 _14172_ ( .A(\u_lsu.pmem[3909] ), .B1(_10231_ ), .B2(_10047_ ), .ZN(_10441_ ) );
AOI21_X1 _14173_ ( .A(fanout_net_14 ), .B1(_10440_ ), .B2(_10441_ ), .ZN(_00352_ ) );
AND2_X2 _14174_ ( .A1(_10423_ ), .A2(_09875_ ), .ZN(_10442_ ) );
BUF_X4 _14175_ ( .A(_10442_ ), .Z(_10443_ ) );
BUF_X4 _14176_ ( .A(_09575_ ), .Z(_10444_ ) );
NAND4_X1 _14177_ ( .A1(_10443_ ), .A2(_10444_ ), .A3(_10385_ ), .A4(_10386_ ), .ZN(_10445_ ) );
BUF_X4 _14178_ ( .A(_09515_ ), .Z(_10446_ ) );
OAI21_X1 _14179_ ( .A(\u_lsu.pmem[7814] ), .B1(_10426_ ), .B2(_10446_ ), .ZN(_10447_ ) );
AOI21_X1 _14180_ ( .A(fanout_net_14 ), .B1(_10445_ ), .B2(_10447_ ), .ZN(_00353_ ) );
BUF_X4 _14181_ ( .A(_09582_ ), .Z(_10448_ ) );
BUF_X4 _14182_ ( .A(_10340_ ), .Z(_10449_ ) );
BUF_X4 _14183_ ( .A(_10033_ ), .Z(_10450_ ) );
NAND4_X1 _14184_ ( .A1(_10443_ ), .A2(_10448_ ), .A3(_10449_ ), .A4(_10450_ ), .ZN(_10451_ ) );
OAI21_X1 _14185_ ( .A(\u_lsu.pmem[7813] ), .B1(_10426_ ), .B2(_10446_ ), .ZN(_10452_ ) );
AOI21_X1 _14186_ ( .A(fanout_net_14 ), .B1(_10451_ ), .B2(_10452_ ), .ZN(_00354_ ) );
BUF_X4 _14187_ ( .A(_08605_ ), .Z(_10453_ ) );
NAND4_X1 _14188_ ( .A1(_10443_ ), .A2(_10453_ ), .A3(_10449_ ), .A4(_10450_ ), .ZN(_10454_ ) );
OAI21_X1 _14189_ ( .A(\u_lsu.pmem[7812] ), .B1(_10426_ ), .B2(_10446_ ), .ZN(_10455_ ) );
AOI21_X1 _14190_ ( .A(fanout_net_14 ), .B1(_10454_ ), .B2(_10455_ ), .ZN(_00355_ ) );
BUF_X4 _14191_ ( .A(_09519_ ), .Z(_10456_ ) );
NAND4_X1 _14192_ ( .A1(_10443_ ), .A2(_10456_ ), .A3(_10449_ ), .A4(_10450_ ), .ZN(_10457_ ) );
OAI21_X1 _14193_ ( .A(\u_lsu.pmem[7811] ), .B1(_10426_ ), .B2(_10446_ ), .ZN(_10458_ ) );
AOI21_X1 _14194_ ( .A(fanout_net_14 ), .B1(_10457_ ), .B2(_10458_ ), .ZN(_00356_ ) );
OAI21_X1 _14195_ ( .A(\u_lsu.pmem[7810] ), .B1(_10426_ ), .B2(_10190_ ), .ZN(_10459_ ) );
NOR3_X1 _14196_ ( .A1(_09533_ ), .A2(_09786_ ), .A3(_09873_ ), .ZN(_10460_ ) );
BUF_X4 _14197_ ( .A(_09950_ ), .Z(_10461_ ) );
NAND4_X1 _14198_ ( .A1(_10460_ ), .A2(_10437_ ), .A3(_10438_ ), .A4(_10461_ ), .ZN(_10462_ ) );
AOI21_X1 _14199_ ( .A(fanout_net_14 ), .B1(_10459_ ), .B2(_10462_ ), .ZN(_00357_ ) );
BUF_X4 _14200_ ( .A(_09543_ ), .Z(_10463_ ) );
NAND4_X1 _14201_ ( .A1(_10443_ ), .A2(_10463_ ), .A3(_10449_ ), .A4(_10450_ ), .ZN(_10464_ ) );
BUF_X4 _14202_ ( .A(_09515_ ), .Z(_10465_ ) );
OAI21_X1 _14203_ ( .A(\u_lsu.pmem[7809] ), .B1(_10426_ ), .B2(_10465_ ), .ZN(_10466_ ) );
AOI21_X1 _14204_ ( .A(fanout_net_14 ), .B1(_10464_ ), .B2(_10466_ ), .ZN(_00358_ ) );
BUF_X4 _14205_ ( .A(_09547_ ), .Z(_10467_ ) );
NAND4_X1 _14206_ ( .A1(_10443_ ), .A2(_10467_ ), .A3(_10449_ ), .A4(_10450_ ), .ZN(_10468_ ) );
OAI21_X1 _14207_ ( .A(\u_lsu.pmem[7808] ), .B1(_10426_ ), .B2(_10465_ ), .ZN(_10469_ ) );
AOI21_X1 _14208_ ( .A(fanout_net_14 ), .B1(_10468_ ), .B2(_10469_ ), .ZN(_00359_ ) );
NAND3_X1 _14209_ ( .A1(_09130_ ), .A2(_10050_ ), .A3(_09556_ ), .ZN(_10470_ ) );
NOR2_X2 _14210_ ( .A1(_09538_ ), .A2(_10470_ ), .ZN(_10471_ ) );
NAND2_X1 _14211_ ( .A1(_10471_ ), .A2(_10326_ ), .ZN(_10472_ ) );
BUF_X4 _14212_ ( .A(_10472_ ), .Z(_10473_ ) );
OAI21_X1 _14213_ ( .A(\u_lsu.pmem[7783] ), .B1(_10360_ ), .B2(_10473_ ), .ZN(_10474_ ) );
BUF_X4 _14214_ ( .A(_10471_ ), .Z(_10475_ ) );
NAND4_X1 _14215_ ( .A1(_10330_ ), .A2(_10366_ ), .A3(_10438_ ), .A4(_10475_ ), .ZN(_10476_ ) );
AOI21_X1 _14216_ ( .A(fanout_net_14 ), .B1(_10474_ ), .B2(_10476_ ), .ZN(_00360_ ) );
OAI21_X1 _14217_ ( .A(\u_lsu.pmem[7782] ), .B1(_10360_ ), .B2(_10473_ ), .ZN(_10477_ ) );
NAND4_X1 _14218_ ( .A1(_09579_ ), .A2(_10366_ ), .A3(_10438_ ), .A4(_10475_ ), .ZN(_10478_ ) );
AOI21_X1 _14219_ ( .A(fanout_net_14 ), .B1(_10477_ ), .B2(_10478_ ), .ZN(_00361_ ) );
OAI21_X1 _14220_ ( .A(\u_lsu.pmem[7781] ), .B1(_10360_ ), .B2(_10473_ ), .ZN(_10479_ ) );
NAND4_X1 _14221_ ( .A1(_09586_ ), .A2(_10366_ ), .A3(_10438_ ), .A4(_10475_ ), .ZN(_10480_ ) );
AOI21_X1 _14222_ ( .A(fanout_net_14 ), .B1(_10479_ ), .B2(_10480_ ), .ZN(_00362_ ) );
NAND4_X1 _14223_ ( .A1(_09736_ ), .A2(_09868_ ), .A3(_09869_ ), .A4(_10450_ ), .ZN(_10481_ ) );
OAI21_X1 _14224_ ( .A(\u_lsu.pmem[4352] ), .B1(_10419_ ), .B2(_09468_ ), .ZN(_10482_ ) );
AOI21_X1 _14225_ ( .A(fanout_net_14 ), .B1(_10481_ ), .B2(_10482_ ), .ZN(_00363_ ) );
OR4_X1 _14226_ ( .A1(_09146_ ), .A2(_10230_ ), .A3(_10113_ ), .A4(_10302_ ), .ZN(_10483_ ) );
OAI21_X1 _14227_ ( .A(\u_lsu.pmem[3908] ), .B1(_10230_ ), .B2(_10047_ ), .ZN(_10484_ ) );
AOI21_X1 _14228_ ( .A(fanout_net_14 ), .B1(_10483_ ), .B2(_10484_ ), .ZN(_00364_ ) );
OAI21_X1 _14229_ ( .A(\u_lsu.pmem[7780] ), .B1(_10360_ ), .B2(_10473_ ), .ZN(_10485_ ) );
BUF_X4 _14230_ ( .A(_09148_ ), .Z(_10486_ ) );
NAND4_X1 _14231_ ( .A1(_10486_ ), .A2(_10366_ ), .A3(_10438_ ), .A4(_10475_ ), .ZN(_10487_ ) );
AOI21_X1 _14232_ ( .A(fanout_net_15 ), .B1(_10485_ ), .B2(_10487_ ), .ZN(_00365_ ) );
OAI21_X1 _14233_ ( .A(\u_lsu.pmem[7779] ), .B1(_10360_ ), .B2(_10473_ ), .ZN(_10488_ ) );
BUF_X4 _14234_ ( .A(_10471_ ), .Z(_10489_ ) );
NAND4_X1 _14235_ ( .A1(_09449_ ), .A2(_10366_ ), .A3(_10438_ ), .A4(_10489_ ), .ZN(_10490_ ) );
AOI21_X1 _14236_ ( .A(fanout_net_15 ), .B1(_10488_ ), .B2(_10490_ ), .ZN(_00366_ ) );
OAI21_X1 _14237_ ( .A(\u_lsu.pmem[7778] ), .B1(_10360_ ), .B2(_10473_ ), .ZN(_10491_ ) );
BUF_X4 _14238_ ( .A(_09611_ ), .Z(_10492_ ) );
NAND4_X1 _14239_ ( .A1(_10492_ ), .A2(_10366_ ), .A3(_10438_ ), .A4(_10489_ ), .ZN(_10493_ ) );
AOI21_X1 _14240_ ( .A(fanout_net_15 ), .B1(_10491_ ), .B2(_10493_ ), .ZN(_00367_ ) );
OAI21_X1 _14241_ ( .A(\u_lsu.pmem[7777] ), .B1(_10360_ ), .B2(_10473_ ), .ZN(_10494_ ) );
NAND4_X1 _14242_ ( .A1(_09698_ ), .A2(_10366_ ), .A3(_10438_ ), .A4(_10489_ ), .ZN(_10495_ ) );
AOI21_X1 _14243_ ( .A(fanout_net_15 ), .B1(_10494_ ), .B2(_10495_ ), .ZN(_00368_ ) );
OAI21_X1 _14244_ ( .A(\u_lsu.pmem[7776] ), .B1(_10360_ ), .B2(_10473_ ), .ZN(_10496_ ) );
NAND4_X1 _14245_ ( .A1(_09622_ ), .A2(_10366_ ), .A3(_10438_ ), .A4(_10489_ ), .ZN(_10497_ ) );
AOI21_X1 _14246_ ( .A(fanout_net_15 ), .B1(_10496_ ), .B2(_10497_ ), .ZN(_00369_ ) );
BUF_X4 _14247_ ( .A(_09572_ ), .Z(_10498_ ) );
AND3_X1 _14248_ ( .A1(_09117_ ), .A2(_09130_ ), .A3(_09947_ ), .ZN(_10499_ ) );
BUF_X4 _14249_ ( .A(_10499_ ), .Z(_10500_ ) );
NAND2_X1 _14250_ ( .A1(_10500_ ), .A2(_10325_ ), .ZN(_10501_ ) );
BUF_X4 _14251_ ( .A(_10501_ ), .Z(_10502_ ) );
OAI21_X1 _14252_ ( .A(\u_lsu.pmem[7751] ), .B1(_10498_ ), .B2(_10502_ ), .ZN(_10503_ ) );
BUF_X4 _14253_ ( .A(_09451_ ), .Z(_10504_ ) );
BUF_X4 _14254_ ( .A(_09878_ ), .Z(_10505_ ) );
BUF_X4 _14255_ ( .A(_10500_ ), .Z(_10506_ ) );
NAND4_X1 _14256_ ( .A1(_10330_ ), .A2(_10504_ ), .A3(_10505_ ), .A4(_10506_ ), .ZN(_10507_ ) );
AOI21_X1 _14257_ ( .A(fanout_net_15 ), .B1(_10503_ ), .B2(_10507_ ), .ZN(_00370_ ) );
OAI21_X1 _14258_ ( .A(\u_lsu.pmem[7750] ), .B1(_10498_ ), .B2(_10502_ ), .ZN(_10508_ ) );
NAND4_X1 _14259_ ( .A1(_09579_ ), .A2(_10504_ ), .A3(_10505_ ), .A4(_10506_ ), .ZN(_10509_ ) );
AOI21_X1 _14260_ ( .A(fanout_net_15 ), .B1(_10508_ ), .B2(_10509_ ), .ZN(_00371_ ) );
OAI21_X1 _14261_ ( .A(\u_lsu.pmem[7749] ), .B1(_10498_ ), .B2(_10502_ ), .ZN(_10510_ ) );
BUF_X4 _14262_ ( .A(_10500_ ), .Z(_10511_ ) );
NAND4_X1 _14263_ ( .A1(_09586_ ), .A2(_10504_ ), .A3(_10505_ ), .A4(_10511_ ), .ZN(_10512_ ) );
AOI21_X1 _14264_ ( .A(fanout_net_15 ), .B1(_10510_ ), .B2(_10512_ ), .ZN(_00372_ ) );
OAI21_X1 _14265_ ( .A(\u_lsu.pmem[7748] ), .B1(_10498_ ), .B2(_10502_ ), .ZN(_10513_ ) );
NAND4_X1 _14266_ ( .A1(_10486_ ), .A2(_10504_ ), .A3(_10505_ ), .A4(_10511_ ), .ZN(_10514_ ) );
AOI21_X1 _14267_ ( .A(fanout_net_15 ), .B1(_10513_ ), .B2(_10514_ ), .ZN(_00373_ ) );
OAI21_X1 _14268_ ( .A(\u_lsu.pmem[7747] ), .B1(_10498_ ), .B2(_10502_ ), .ZN(_10515_ ) );
NAND4_X1 _14269_ ( .A1(_09449_ ), .A2(_10504_ ), .A3(_10505_ ), .A4(_10511_ ), .ZN(_10516_ ) );
AOI21_X1 _14270_ ( .A(fanout_net_15 ), .B1(_10515_ ), .B2(_10516_ ), .ZN(_00374_ ) );
OR4_X1 _14271_ ( .A1(_09969_ ), .A2(_10230_ ), .A3(_10113_ ), .A4(_10302_ ), .ZN(_10517_ ) );
BUF_X4 _14272_ ( .A(_10046_ ), .Z(_10518_ ) );
OAI21_X1 _14273_ ( .A(\u_lsu.pmem[3907] ), .B1(_10230_ ), .B2(_10518_ ), .ZN(_10519_ ) );
AOI21_X1 _14274_ ( .A(fanout_net_15 ), .B1(_10517_ ), .B2(_10519_ ), .ZN(_00375_ ) );
OAI21_X1 _14275_ ( .A(\u_lsu.pmem[7746] ), .B1(_10498_ ), .B2(_10502_ ), .ZN(_10520_ ) );
NAND4_X1 _14276_ ( .A1(_10492_ ), .A2(_10504_ ), .A3(_10505_ ), .A4(_10511_ ), .ZN(_10521_ ) );
AOI21_X1 _14277_ ( .A(fanout_net_15 ), .B1(_10520_ ), .B2(_10521_ ), .ZN(_00376_ ) );
OAI21_X1 _14278_ ( .A(\u_lsu.pmem[7745] ), .B1(_10498_ ), .B2(_10502_ ), .ZN(_10522_ ) );
NAND4_X1 _14279_ ( .A1(_09698_ ), .A2(_10504_ ), .A3(_10505_ ), .A4(_10511_ ), .ZN(_10523_ ) );
AOI21_X1 _14280_ ( .A(fanout_net_15 ), .B1(_10522_ ), .B2(_10523_ ), .ZN(_00377_ ) );
OAI21_X1 _14281_ ( .A(\u_lsu.pmem[7744] ), .B1(_10498_ ), .B2(_10502_ ), .ZN(_10524_ ) );
BUF_X4 _14282_ ( .A(_09621_ ), .Z(_10525_ ) );
NAND4_X1 _14283_ ( .A1(_10525_ ), .A2(_10504_ ), .A3(_10505_ ), .A4(_10511_ ), .ZN(_10526_ ) );
AOI21_X1 _14284_ ( .A(fanout_net_15 ), .B1(_10524_ ), .B2(_10526_ ), .ZN(_00378_ ) );
AND3_X2 _14285_ ( .A1(_09663_ ), .A2(_09760_ ), .A3(_09762_ ), .ZN(_10527_ ) );
NAND4_X1 _14286_ ( .A1(_10527_ ), .A2(_10395_ ), .A3(_10449_ ), .A4(_10450_ ), .ZN(_10528_ ) );
BUF_X4 _14287_ ( .A(_09482_ ), .Z(_10529_ ) );
NOR3_X1 _14288_ ( .A1(_09129_ ), .A2(_10529_ ), .A3(_09126_ ), .ZN(_10530_ ) );
AND2_X2 _14289_ ( .A1(_10530_ ), .A2(_09743_ ), .ZN(_10531_ ) );
NAND2_X2 _14290_ ( .A1(_10531_ ), .A2(_09877_ ), .ZN(_10532_ ) );
BUF_X4 _14291_ ( .A(_10532_ ), .Z(_10533_ ) );
OAI21_X1 _14292_ ( .A(\u_lsu.pmem[7719] ), .B1(_10419_ ), .B2(_10533_ ), .ZN(_10534_ ) );
AOI21_X1 _14293_ ( .A(fanout_net_15 ), .B1(_10528_ ), .B2(_10534_ ), .ZN(_00379_ ) );
AND3_X2 _14294_ ( .A1(_09680_ ), .A2(_09760_ ), .A3(_09762_ ), .ZN(_10535_ ) );
NAND4_X1 _14295_ ( .A1(_10535_ ), .A2(_10395_ ), .A3(_10449_ ), .A4(_10450_ ), .ZN(_10536_ ) );
OAI21_X1 _14296_ ( .A(\u_lsu.pmem[7718] ), .B1(_10419_ ), .B2(_10533_ ), .ZN(_10537_ ) );
AOI21_X1 _14297_ ( .A(fanout_net_15 ), .B1(_10536_ ), .B2(_10537_ ), .ZN(_00380_ ) );
AND3_X2 _14298_ ( .A1(_09684_ ), .A2(_09760_ ), .A3(_09762_ ), .ZN(_10538_ ) );
NAND4_X1 _14299_ ( .A1(_10538_ ), .A2(_10395_ ), .A3(_10449_ ), .A4(_10450_ ), .ZN(_10539_ ) );
OAI21_X1 _14300_ ( .A(\u_lsu.pmem[7717] ), .B1(_10419_ ), .B2(_10533_ ), .ZN(_10540_ ) );
AOI21_X1 _14301_ ( .A(fanout_net_15 ), .B1(_10539_ ), .B2(_10540_ ), .ZN(_00381_ ) );
OAI21_X1 _14302_ ( .A(\u_lsu.pmem[7716] ), .B1(_10498_ ), .B2(_10533_ ), .ZN(_10541_ ) );
BUF_X4 _14303_ ( .A(_10531_ ), .Z(_10542_ ) );
NAND4_X1 _14304_ ( .A1(_10486_ ), .A2(_10504_ ), .A3(_10505_ ), .A4(_10542_ ), .ZN(_10543_ ) );
AOI21_X1 _14305_ ( .A(fanout_net_15 ), .B1(_10541_ ), .B2(_10543_ ), .ZN(_00382_ ) );
OAI21_X1 _14306_ ( .A(\u_lsu.pmem[7715] ), .B1(_10498_ ), .B2(_10533_ ), .ZN(_10544_ ) );
NAND4_X1 _14307_ ( .A1(_09449_ ), .A2(_10504_ ), .A3(_10505_ ), .A4(_10542_ ), .ZN(_10545_ ) );
AOI21_X1 _14308_ ( .A(fanout_net_15 ), .B1(_10544_ ), .B2(_10545_ ), .ZN(_00383_ ) );
BUF_X4 _14309_ ( .A(_09572_ ), .Z(_10546_ ) );
OAI21_X1 _14310_ ( .A(\u_lsu.pmem[7714] ), .B1(_10546_ ), .B2(_10533_ ), .ZN(_10547_ ) );
BUF_X8 _14311_ ( .A(_09450_ ), .Z(_10548_ ) );
BUF_X4 _14312_ ( .A(_10548_ ), .Z(_10549_ ) );
BUF_X4 _14313_ ( .A(_09878_ ), .Z(_10550_ ) );
NAND4_X1 _14314_ ( .A1(_10492_ ), .A2(_10549_ ), .A3(_10550_ ), .A4(_10542_ ), .ZN(_10551_ ) );
AOI21_X1 _14315_ ( .A(fanout_net_15 ), .B1(_10547_ ), .B2(_10551_ ), .ZN(_00384_ ) );
OAI21_X1 _14316_ ( .A(\u_lsu.pmem[7713] ), .B1(_10546_ ), .B2(_10533_ ), .ZN(_10552_ ) );
NAND4_X1 _14317_ ( .A1(_09698_ ), .A2(_10549_ ), .A3(_10550_ ), .A4(_10542_ ), .ZN(_10553_ ) );
AOI21_X1 _14318_ ( .A(fanout_net_15 ), .B1(_10552_ ), .B2(_10553_ ), .ZN(_00385_ ) );
OR4_X1 _14319_ ( .A1(_09973_ ), .A2(_10229_ ), .A3(_10045_ ), .A4(_10302_ ), .ZN(_10554_ ) );
OAI21_X1 _14320_ ( .A(\u_lsu.pmem[3906] ), .B1(_10230_ ), .B2(_10518_ ), .ZN(_10555_ ) );
AOI21_X1 _14321_ ( .A(fanout_net_15 ), .B1(_10554_ ), .B2(_10555_ ), .ZN(_00386_ ) );
NOR3_X4 _14322_ ( .A1(_09701_ ), .A2(_09669_ ), .A3(_09873_ ), .ZN(_10556_ ) );
BUF_X4 _14323_ ( .A(_10126_ ), .Z(_10557_ ) );
NAND4_X1 _14324_ ( .A1(_10556_ ), .A2(_10557_ ), .A3(_10449_ ), .A4(_10450_ ), .ZN(_10558_ ) );
OAI21_X1 _14325_ ( .A(\u_lsu.pmem[7712] ), .B1(_10419_ ), .B2(_10533_ ), .ZN(_10559_ ) );
AOI21_X1 _14326_ ( .A(fanout_net_15 ), .B1(_10558_ ), .B2(_10559_ ), .ZN(_00387_ ) );
AND2_X1 _14327_ ( .A1(_09114_ ), .A2(_10252_ ), .ZN(_10560_ ) );
AND2_X1 _14328_ ( .A1(_10560_ ), .A2(_09489_ ), .ZN(_10561_ ) );
AND2_X1 _14329_ ( .A1(_10561_ ), .A2(_09491_ ), .ZN(_10562_ ) );
INV_X1 _14330_ ( .A(_10562_ ), .ZN(_10563_ ) );
BUF_X4 _14331_ ( .A(_10563_ ), .Z(_10564_ ) );
OAI21_X1 _14332_ ( .A(\u_lsu.pmem[7687] ), .B1(_10564_ ), .B2(_10240_ ), .ZN(_10565_ ) );
BUF_X4 _14333_ ( .A(_10561_ ), .Z(_10566_ ) );
NAND4_X1 _14334_ ( .A1(_10566_ ), .A2(_09603_ ), .A3(_10244_ ), .A4(_10273_ ), .ZN(_10567_ ) );
AOI21_X1 _14335_ ( .A(fanout_net_15 ), .B1(_10565_ ), .B2(_10567_ ), .ZN(_00388_ ) );
OAI21_X1 _14336_ ( .A(\u_lsu.pmem[7686] ), .B1(_10564_ ), .B2(_10240_ ), .ZN(_10568_ ) );
NAND4_X1 _14337_ ( .A1(_10566_ ), .A2(_10185_ ), .A3(_10244_ ), .A4(_10273_ ), .ZN(_10569_ ) );
AOI21_X1 _14338_ ( .A(fanout_net_15 ), .B1(_10568_ ), .B2(_10569_ ), .ZN(_00389_ ) );
OAI21_X1 _14339_ ( .A(\u_lsu.pmem[7685] ), .B1(_10564_ ), .B2(_10240_ ), .ZN(_10570_ ) );
NAND4_X1 _14340_ ( .A1(_10566_ ), .A2(_10188_ ), .A3(_10244_ ), .A4(_10273_ ), .ZN(_10571_ ) );
AOI21_X1 _14341_ ( .A(fanout_net_15 ), .B1(_10570_ ), .B2(_10571_ ), .ZN(_00390_ ) );
BUF_X4 _14342_ ( .A(_10070_ ), .Z(_10572_ ) );
OAI21_X1 _14343_ ( .A(\u_lsu.pmem[7684] ), .B1(_10564_ ), .B2(_10572_ ), .ZN(_10573_ ) );
NAND4_X1 _14344_ ( .A1(_10566_ ), .A2(_10192_ ), .A3(_10244_ ), .A4(_10273_ ), .ZN(_10574_ ) );
AOI21_X1 _14345_ ( .A(fanout_net_15 ), .B1(_10573_ ), .B2(_10574_ ), .ZN(_00391_ ) );
AND2_X2 _14346_ ( .A1(_09448_ ), .A2(_10560_ ), .ZN(_10575_ ) );
BUF_X4 _14347_ ( .A(_10046_ ), .Z(_10576_ ) );
BUF_X4 _14348_ ( .A(_10287_ ), .Z(_10577_ ) );
BUF_X8 _14349_ ( .A(_09877_ ), .Z(_10578_ ) );
BUF_X4 _14350_ ( .A(_10578_ ), .Z(_10579_ ) );
NAND4_X1 _14351_ ( .A1(_10575_ ), .A2(_10576_ ), .A3(_10577_ ), .A4(_10579_ ), .ZN(_10580_ ) );
OAI21_X1 _14352_ ( .A(\u_lsu.pmem[7683] ), .B1(_10563_ ), .B2(_10140_ ), .ZN(_10581_ ) );
AOI21_X1 _14353_ ( .A(fanout_net_15 ), .B1(_10580_ ), .B2(_10581_ ), .ZN(_00392_ ) );
NOR2_X1 _14354_ ( .A1(_09145_ ), .A2(_09464_ ), .ZN(_10582_ ) );
NAND3_X1 _14355_ ( .A1(_10582_ ), .A2(_09474_ ), .A3(_09669_ ), .ZN(_10583_ ) );
NOR2_X1 _14356_ ( .A1(_10583_ ), .A2(_09774_ ), .ZN(_10584_ ) );
BUF_X2 _14357_ ( .A(_09605_ ), .Z(\alu_result_out[8] ) );
BUF_X4 _14358_ ( .A(_10287_ ), .Z(_10585_ ) );
NAND4_X1 _14359_ ( .A1(_10584_ ), .A2(_10576_ ), .A3(\alu_result_out[8] ), .A4(_10585_ ), .ZN(_10586_ ) );
OAI21_X1 _14360_ ( .A(\u_lsu.pmem[7682] ), .B1(_10563_ ), .B2(_10140_ ), .ZN(_10587_ ) );
AOI21_X1 _14361_ ( .A(fanout_net_15 ), .B1(_10586_ ), .B2(_10587_ ), .ZN(_00393_ ) );
OAI21_X1 _14362_ ( .A(\u_lsu.pmem[7681] ), .B1(_10564_ ), .B2(_10572_ ), .ZN(_10588_ ) );
BUF_X4 _14363_ ( .A(_10041_ ), .Z(_10589_ ) );
NAND4_X1 _14364_ ( .A1(_10566_ ), .A2(_09923_ ), .A3(_10589_ ), .A4(_10273_ ), .ZN(_10590_ ) );
AOI21_X1 _14365_ ( .A(fanout_net_15 ), .B1(_10588_ ), .B2(_10590_ ), .ZN(_00394_ ) );
AND2_X2 _14366_ ( .A1(_09620_ ), .A2(_10560_ ), .ZN(_10591_ ) );
BUF_X8 _14367_ ( .A(_09471_ ), .Z(_10592_ ) );
BUF_X4 _14368_ ( .A(_10592_ ), .Z(_10593_ ) );
NAND4_X1 _14369_ ( .A1(_10591_ ), .A2(_10557_ ), .A3(_10449_ ), .A4(_10593_ ), .ZN(_10594_ ) );
OAI21_X1 _14370_ ( .A(\u_lsu.pmem[7680] ), .B1(_10563_ ), .B2(_10140_ ), .ZN(_10595_ ) );
AOI21_X1 _14371_ ( .A(fanout_net_16 ), .B1(_10594_ ), .B2(_10595_ ), .ZN(_00395_ ) );
AND3_X1 _14372_ ( .A1(_10397_ ), .A2(_09505_ ), .A3(_10052_ ), .ZN(_10596_ ) );
NAND2_X4 _14373_ ( .A1(_10596_ ), .A2(_10326_ ), .ZN(_10597_ ) );
BUF_X4 _14374_ ( .A(_10597_ ), .Z(_10598_ ) );
OAI21_X1 _14375_ ( .A(\u_lsu.pmem[7655] ), .B1(_10546_ ), .B2(_10598_ ), .ZN(_10599_ ) );
NAND4_X1 _14376_ ( .A1(_10330_ ), .A2(_10549_ ), .A3(_10550_ ), .A4(_10596_ ), .ZN(_10600_ ) );
AOI21_X1 _14377_ ( .A(fanout_net_16 ), .B1(_10599_ ), .B2(_10600_ ), .ZN(_00396_ ) );
OR4_X1 _14378_ ( .A1(_09977_ ), .A2(_10229_ ), .A3(_10045_ ), .A4(_10302_ ), .ZN(_10601_ ) );
OAI21_X1 _14379_ ( .A(\u_lsu.pmem[3905] ), .B1(_10230_ ), .B2(_10518_ ), .ZN(_10602_ ) );
AOI21_X1 _14380_ ( .A(fanout_net_16 ), .B1(_10601_ ), .B2(_10602_ ), .ZN(_00397_ ) );
NOR2_X1 _14381_ ( .A1(_10060_ ), .A2(_09536_ ), .ZN(_10603_ ) );
BUF_X4 _14382_ ( .A(_10340_ ), .Z(_10604_ ) );
NAND4_X1 _14383_ ( .A1(_10603_ ), .A2(_10557_ ), .A3(_10604_ ), .A4(_10593_ ), .ZN(_10605_ ) );
OAI21_X1 _14384_ ( .A(\u_lsu.pmem[7654] ), .B1(_10419_ ), .B2(_10598_ ), .ZN(_10606_ ) );
AOI21_X1 _14385_ ( .A(fanout_net_16 ), .B1(_10605_ ), .B2(_10606_ ), .ZN(_00398_ ) );
BUF_X4 _14386_ ( .A(_10093_ ), .Z(_10607_ ) );
AND2_X2 _14387_ ( .A1(_10073_ ), .A2(_10607_ ), .ZN(_10608_ ) );
NAND4_X1 _14388_ ( .A1(_10608_ ), .A2(_10576_ ), .A3(_10577_ ), .A4(_10579_ ), .ZN(_10609_ ) );
OAI21_X1 _14389_ ( .A(\u_lsu.pmem[7653] ), .B1(_10419_ ), .B2(_10598_ ), .ZN(_10610_ ) );
AOI21_X1 _14390_ ( .A(fanout_net_16 ), .B1(_10609_ ), .B2(_10610_ ), .ZN(_00399_ ) );
AND2_X4 _14391_ ( .A1(_10078_ ), .A2(_10607_ ), .ZN(_10611_ ) );
NAND4_X1 _14392_ ( .A1(_10611_ ), .A2(_10576_ ), .A3(_10577_ ), .A4(_10579_ ), .ZN(_10612_ ) );
OAI21_X1 _14393_ ( .A(\u_lsu.pmem[7652] ), .B1(_10419_ ), .B2(_10598_ ), .ZN(_10613_ ) );
AOI21_X1 _14394_ ( .A(fanout_net_16 ), .B1(_10612_ ), .B2(_10613_ ), .ZN(_00400_ ) );
AND2_X2 _14395_ ( .A1(_10083_ ), .A2(_10607_ ), .ZN(_10614_ ) );
NAND4_X1 _14396_ ( .A1(_10614_ ), .A2(_10576_ ), .A3(_10577_ ), .A4(_10579_ ), .ZN(_10615_ ) );
OAI21_X1 _14397_ ( .A(\u_lsu.pmem[7651] ), .B1(_10419_ ), .B2(_10598_ ), .ZN(_10616_ ) );
AOI21_X1 _14398_ ( .A(fanout_net_16 ), .B1(_10615_ ), .B2(_10616_ ), .ZN(_00401_ ) );
AND2_X2 _14399_ ( .A1(_10087_ ), .A2(_10607_ ), .ZN(_10617_ ) );
NAND4_X1 _14400_ ( .A1(_10617_ ), .A2(_10576_ ), .A3(_10577_ ), .A4(_10579_ ), .ZN(_10618_ ) );
BUF_X4 _14401_ ( .A(_10036_ ), .Z(_10619_ ) );
OAI21_X1 _14402_ ( .A(\u_lsu.pmem[7650] ), .B1(_10619_ ), .B2(_10598_ ), .ZN(_10620_ ) );
AOI21_X1 _14403_ ( .A(fanout_net_16 ), .B1(_10618_ ), .B2(_10620_ ), .ZN(_00402_ ) );
NOR3_X4 _14404_ ( .A1(_09783_ ), .A2(_09535_ ), .A3(_09536_ ), .ZN(_10621_ ) );
NAND4_X1 _14405_ ( .A1(_10621_ ), .A2(_10557_ ), .A3(_10604_ ), .A4(_10593_ ), .ZN(_10622_ ) );
OAI21_X1 _14406_ ( .A(\u_lsu.pmem[7649] ), .B1(_10619_ ), .B2(_10598_ ), .ZN(_10623_ ) );
AOI21_X1 _14407_ ( .A(fanout_net_16 ), .B1(_10622_ ), .B2(_10623_ ), .ZN(_00403_ ) );
AND2_X2 _14408_ ( .A1(_10097_ ), .A2(_10607_ ), .ZN(_10624_ ) );
NAND4_X1 _14409_ ( .A1(_10624_ ), .A2(\alu_result_out[7] ), .A3(_10604_ ), .A4(_10593_ ), .ZN(_10625_ ) );
OAI21_X1 _14410_ ( .A(\u_lsu.pmem[7648] ), .B1(_10619_ ), .B2(_10598_ ), .ZN(_10626_ ) );
AOI21_X1 _14411_ ( .A(fanout_net_16 ), .B1(_10625_ ), .B2(_10626_ ), .ZN(_00404_ ) );
AND3_X1 _14412_ ( .A1(_09118_ ), .A2(_09505_ ), .A3(_10102_ ), .ZN(_10627_ ) );
NAND2_X4 _14413_ ( .A1(_10627_ ), .A2(_10326_ ), .ZN(_10628_ ) );
BUF_X4 _14414_ ( .A(_10628_ ), .Z(_10629_ ) );
OAI21_X1 _14415_ ( .A(\u_lsu.pmem[7623] ), .B1(_10546_ ), .B2(_10629_ ), .ZN(_10630_ ) );
NAND4_X1 _14416_ ( .A1(_10330_ ), .A2(_10549_ ), .A3(_10550_ ), .A4(_10627_ ), .ZN(_10631_ ) );
AOI21_X1 _14417_ ( .A(fanout_net_16 ), .B1(_10630_ ), .B2(_10631_ ), .ZN(_00405_ ) );
AND2_X2 _14418_ ( .A1(_10116_ ), .A2(_10607_ ), .ZN(_10632_ ) );
NAND4_X1 _14419_ ( .A1(_10632_ ), .A2(_10576_ ), .A3(_10577_ ), .A4(_10579_ ), .ZN(_10633_ ) );
OAI21_X1 _14420_ ( .A(\u_lsu.pmem[7622] ), .B1(_10619_ ), .B2(_10629_ ), .ZN(_10634_ ) );
AOI21_X1 _14421_ ( .A(fanout_net_16 ), .B1(_10633_ ), .B2(_10634_ ), .ZN(_00406_ ) );
AND2_X2 _14422_ ( .A1(_10120_ ), .A2(_10607_ ), .ZN(_10635_ ) );
BUF_X4 _14423_ ( .A(_10046_ ), .Z(_10636_ ) );
NAND4_X1 _14424_ ( .A1(_10635_ ), .A2(_10636_ ), .A3(_10577_ ), .A4(_10579_ ), .ZN(_10637_ ) );
OAI21_X1 _14425_ ( .A(\u_lsu.pmem[7621] ), .B1(_10619_ ), .B2(_10629_ ), .ZN(_10638_ ) );
AOI21_X1 _14426_ ( .A(fanout_net_16 ), .B1(_10637_ ), .B2(_10638_ ), .ZN(_00407_ ) );
OR4_X1 _14427_ ( .A1(_09497_ ), .A2(_10229_ ), .A3(_10045_ ), .A4(_10302_ ), .ZN(_10639_ ) );
OAI21_X1 _14428_ ( .A(\u_lsu.pmem[3904] ), .B1(_10230_ ), .B2(_10518_ ), .ZN(_10640_ ) );
AOI21_X1 _14429_ ( .A(fanout_net_16 ), .B1(_10639_ ), .B2(_10640_ ), .ZN(_00408_ ) );
AND2_X2 _14430_ ( .A1(_10124_ ), .A2(_10607_ ), .ZN(_10641_ ) );
BUF_X4 _14431_ ( .A(_10287_ ), .Z(_10642_ ) );
NAND4_X1 _14432_ ( .A1(_10641_ ), .A2(_10636_ ), .A3(_10642_ ), .A4(_10579_ ), .ZN(_10643_ ) );
OAI21_X1 _14433_ ( .A(\u_lsu.pmem[7620] ), .B1(_10619_ ), .B2(_10629_ ), .ZN(_10644_ ) );
AOI21_X1 _14434_ ( .A(fanout_net_16 ), .B1(_10643_ ), .B2(_10644_ ), .ZN(_00409_ ) );
AND2_X2 _14435_ ( .A1(_10130_ ), .A2(_10607_ ), .ZN(_10645_ ) );
BUF_X4 _14436_ ( .A(_10578_ ), .Z(_10646_ ) );
NAND4_X1 _14437_ ( .A1(_10645_ ), .A2(_10636_ ), .A3(_10642_ ), .A4(_10646_ ), .ZN(_10647_ ) );
OAI21_X1 _14438_ ( .A(\u_lsu.pmem[7619] ), .B1(_10619_ ), .B2(_10629_ ), .ZN(_10648_ ) );
AOI21_X1 _14439_ ( .A(fanout_net_16 ), .B1(_10647_ ), .B2(_10648_ ), .ZN(_00410_ ) );
AND2_X2 _14440_ ( .A1(_10134_ ), .A2(_10607_ ), .ZN(_10649_ ) );
NAND4_X1 _14441_ ( .A1(_10649_ ), .A2(_10636_ ), .A3(_10642_ ), .A4(_10646_ ), .ZN(_10650_ ) );
OAI21_X1 _14442_ ( .A(\u_lsu.pmem[7618] ), .B1(_10619_ ), .B2(_10629_ ), .ZN(_10651_ ) );
AOI21_X1 _14443_ ( .A(fanout_net_16 ), .B1(_10650_ ), .B2(_10651_ ), .ZN(_00411_ ) );
NOR3_X4 _14444_ ( .A1(_09830_ ), .A2(_09535_ ), .A3(_09536_ ), .ZN(_10652_ ) );
NAND4_X1 _14445_ ( .A1(_10652_ ), .A2(_10557_ ), .A3(_10604_ ), .A4(_10593_ ), .ZN(_10653_ ) );
OAI21_X1 _14446_ ( .A(\u_lsu.pmem[7617] ), .B1(_10619_ ), .B2(_10629_ ), .ZN(_10654_ ) );
AOI21_X1 _14447_ ( .A(fanout_net_16 ), .B1(_10653_ ), .B2(_10654_ ), .ZN(_00412_ ) );
AND2_X2 _14448_ ( .A1(_10142_ ), .A2(_09986_ ), .ZN(_10655_ ) );
NAND4_X1 _14449_ ( .A1(_10655_ ), .A2(_10636_ ), .A3(_10642_ ), .A4(_10646_ ), .ZN(_10656_ ) );
OAI21_X1 _14450_ ( .A(\u_lsu.pmem[7616] ), .B1(_10619_ ), .B2(_10629_ ), .ZN(_10657_ ) );
AOI21_X1 _14451_ ( .A(fanout_net_16 ), .B1(_10656_ ), .B2(_10657_ ), .ZN(_00413_ ) );
AND2_X2 _14452_ ( .A1(_10147_ ), .A2(_09986_ ), .ZN(_10658_ ) );
NAND4_X1 _14453_ ( .A1(_10658_ ), .A2(\alu_result_out[7] ), .A3(_10604_ ), .A4(_10593_ ), .ZN(_10659_ ) );
BUF_X4 _14454_ ( .A(_10036_ ), .Z(_10660_ ) );
AND3_X2 _14455_ ( .A1(_10397_ ), .A2(_09505_ ), .A3(_10165_ ), .ZN(_10661_ ) );
NAND2_X1 _14456_ ( .A1(_10661_ ), .A2(_10326_ ), .ZN(_10662_ ) );
BUF_X4 _14457_ ( .A(_10662_ ), .Z(_10663_ ) );
OAI21_X1 _14458_ ( .A(\u_lsu.pmem[7591] ), .B1(_10660_ ), .B2(_10663_ ), .ZN(_10664_ ) );
AOI21_X1 _14459_ ( .A(fanout_net_16 ), .B1(_10659_ ), .B2(_10664_ ), .ZN(_00414_ ) );
NOR2_X1 _14460_ ( .A1(_10155_ ), .A2(_09536_ ), .ZN(_10665_ ) );
NAND4_X1 _14461_ ( .A1(_10665_ ), .A2(_10557_ ), .A3(_10604_ ), .A4(_10593_ ), .ZN(_10666_ ) );
OAI21_X1 _14462_ ( .A(\u_lsu.pmem[7590] ), .B1(_10660_ ), .B2(_10663_ ), .ZN(_10667_ ) );
AOI21_X1 _14463_ ( .A(fanout_net_16 ), .B1(_10666_ ), .B2(_10667_ ), .ZN(_00415_ ) );
AND2_X2 _14464_ ( .A1(_10159_ ), .A2(_09986_ ), .ZN(_10668_ ) );
NAND4_X1 _14465_ ( .A1(_10668_ ), .A2(_10636_ ), .A3(_10642_ ), .A4(_10646_ ), .ZN(_10669_ ) );
OAI21_X1 _14466_ ( .A(\u_lsu.pmem[7589] ), .B1(_10660_ ), .B2(_10663_ ), .ZN(_10670_ ) );
AOI21_X1 _14467_ ( .A(fanout_net_16 ), .B1(_10669_ ), .B2(_10670_ ), .ZN(_00416_ ) );
AND3_X2 _14468_ ( .A1(_09148_ ), .A2(_09986_ ), .A3(_10165_ ), .ZN(_10671_ ) );
NAND4_X1 _14469_ ( .A1(_10671_ ), .A2(_10557_ ), .A3(_10604_ ), .A4(_10593_ ), .ZN(_10672_ ) );
OAI21_X1 _14470_ ( .A(\u_lsu.pmem[7588] ), .B1(_10660_ ), .B2(_10663_ ), .ZN(_10673_ ) );
AOI21_X1 _14471_ ( .A(fanout_net_16 ), .B1(_10672_ ), .B2(_10673_ ), .ZN(_00417_ ) );
AND3_X2 _14472_ ( .A1(_09447_ ), .A2(_09986_ ), .A3(_10165_ ), .ZN(_10674_ ) );
NAND4_X1 _14473_ ( .A1(_10674_ ), .A2(_10557_ ), .A3(_10604_ ), .A4(_10593_ ), .ZN(_10675_ ) );
OAI21_X1 _14474_ ( .A(\u_lsu.pmem[7587] ), .B1(_10660_ ), .B2(_10663_ ), .ZN(_10676_ ) );
AOI21_X1 _14475_ ( .A(fanout_net_16 ), .B1(_10675_ ), .B2(_10676_ ), .ZN(_00418_ ) );
NAND4_X1 _14476_ ( .A1(_10250_ ), .A2(_10557_ ), .A3(_10604_ ), .A4(_09998_ ), .ZN(_10677_ ) );
OAI21_X1 _14477_ ( .A(\u_lsu.pmem[3879] ), .B1(_10257_ ), .B2(_10518_ ), .ZN(_10678_ ) );
AOI21_X1 _14478_ ( .A(fanout_net_16 ), .B1(_10677_ ), .B2(_10678_ ), .ZN(_00419_ ) );
AND3_X2 _14479_ ( .A1(_09611_ ), .A2(_09986_ ), .A3(_10165_ ), .ZN(_10679_ ) );
NAND4_X1 _14480_ ( .A1(_10679_ ), .A2(_10557_ ), .A3(_10604_ ), .A4(_10593_ ), .ZN(_10680_ ) );
OAI21_X1 _14481_ ( .A(\u_lsu.pmem[7586] ), .B1(_10660_ ), .B2(_10663_ ), .ZN(_10681_ ) );
AOI21_X1 _14482_ ( .A(fanout_net_16 ), .B1(_10680_ ), .B2(_10681_ ), .ZN(_00420_ ) );
AND3_X2 _14483_ ( .A1(_09615_ ), .A2(_09986_ ), .A3(_10165_ ), .ZN(_10682_ ) );
BUF_X4 _14484_ ( .A(_10126_ ), .Z(_10683_ ) );
BUF_X4 _14485_ ( .A(_10340_ ), .Z(_10684_ ) );
BUF_X4 _14486_ ( .A(_10592_ ), .Z(_10685_ ) );
NAND4_X1 _14487_ ( .A1(_10682_ ), .A2(_10683_ ), .A3(_10684_ ), .A4(_10685_ ), .ZN(_10686_ ) );
OAI21_X1 _14488_ ( .A(\u_lsu.pmem[7585] ), .B1(_10660_ ), .B2(_10663_ ), .ZN(_10687_ ) );
AOI21_X1 _14489_ ( .A(fanout_net_16 ), .B1(_10686_ ), .B2(_10687_ ), .ZN(_00421_ ) );
OAI21_X1 _14490_ ( .A(\u_lsu.pmem[7584] ), .B1(_10546_ ), .B2(_10663_ ), .ZN(_10688_ ) );
NAND4_X1 _14491_ ( .A1(_10525_ ), .A2(_10549_ ), .A3(_10550_ ), .A4(_10661_ ), .ZN(_10689_ ) );
AOI21_X1 _14492_ ( .A(fanout_net_16 ), .B1(_10688_ ), .B2(_10689_ ), .ZN(_00422_ ) );
AND3_X1 _14493_ ( .A1(_09504_ ), .A2(_09505_ ), .A3(_10397_ ), .ZN(_10690_ ) );
NAND2_X1 _14494_ ( .A1(_10690_ ), .A2(_09877_ ), .ZN(_10691_ ) );
BUF_X4 _14495_ ( .A(_10691_ ), .Z(_10692_ ) );
OAI21_X1 _14496_ ( .A(\u_lsu.pmem[7559] ), .B1(_10692_ ), .B2(_10190_ ), .ZN(_10693_ ) );
BUF_X4 _14497_ ( .A(_10690_ ), .Z(_10694_ ) );
BUF_X4 _14498_ ( .A(_10694_ ), .Z(_10695_ ) );
NAND4_X1 _14499_ ( .A1(_10695_ ), .A2(_09603_ ), .A3(_10550_ ), .A4(_10461_ ), .ZN(_10696_ ) );
AOI21_X1 _14500_ ( .A(fanout_net_16 ), .B1(_10693_ ), .B2(_10696_ ), .ZN(_00423_ ) );
OAI21_X1 _14501_ ( .A(\u_lsu.pmem[7558] ), .B1(_10692_ ), .B2(_10190_ ), .ZN(_10697_ ) );
NAND4_X1 _14502_ ( .A1(_10695_ ), .A2(_10185_ ), .A3(_10550_ ), .A4(_10461_ ), .ZN(_10698_ ) );
AOI21_X1 _14503_ ( .A(fanout_net_16 ), .B1(_10697_ ), .B2(_10698_ ), .ZN(_00424_ ) );
OAI21_X1 _14504_ ( .A(\u_lsu.pmem[7557] ), .B1(_10692_ ), .B2(_10190_ ), .ZN(_10699_ ) );
NAND4_X1 _14505_ ( .A1(_10695_ ), .A2(_10188_ ), .A3(_10550_ ), .A4(_10461_ ), .ZN(_10700_ ) );
AOI21_X1 _14506_ ( .A(fanout_net_17 ), .B1(_10699_ ), .B2(_10700_ ), .ZN(_00425_ ) );
BUF_X4 _14507_ ( .A(_09443_ ), .Z(_10701_ ) );
OAI21_X1 _14508_ ( .A(\u_lsu.pmem[7556] ), .B1(_10692_ ), .B2(_10701_ ), .ZN(_10702_ ) );
NAND4_X1 _14509_ ( .A1(_10695_ ), .A2(_10192_ ), .A3(_10550_ ), .A4(_10461_ ), .ZN(_10703_ ) );
AOI21_X1 _14510_ ( .A(fanout_net_17 ), .B1(_10702_ ), .B2(_10703_ ), .ZN(_00426_ ) );
OAI21_X1 _14511_ ( .A(\u_lsu.pmem[7555] ), .B1(_10692_ ), .B2(_10701_ ), .ZN(_10704_ ) );
NAND4_X1 _14512_ ( .A1(_10695_ ), .A2(_09520_ ), .A3(_10550_ ), .A4(_10461_ ), .ZN(_10705_ ) );
AOI21_X1 _14513_ ( .A(fanout_net_17 ), .B1(_10704_ ), .B2(_10705_ ), .ZN(_00427_ ) );
OAI21_X1 _14514_ ( .A(\u_lsu.pmem[7554] ), .B1(_10692_ ), .B2(_10701_ ), .ZN(_10706_ ) );
BUF_X4 _14515_ ( .A(_09878_ ), .Z(_10707_ ) );
NAND4_X1 _14516_ ( .A1(_09537_ ), .A2(_10437_ ), .A3(_10707_ ), .A4(_10461_ ), .ZN(_10708_ ) );
AOI21_X1 _14517_ ( .A(fanout_net_17 ), .B1(_10706_ ), .B2(_10708_ ), .ZN(_00428_ ) );
OAI21_X1 _14518_ ( .A(\u_lsu.pmem[7553] ), .B1(_10692_ ), .B2(_10701_ ), .ZN(_10709_ ) );
NAND4_X1 _14519_ ( .A1(_10695_ ), .A2(_09923_ ), .A3(_10707_ ), .A4(_10461_ ), .ZN(_10710_ ) );
AOI21_X1 _14520_ ( .A(fanout_net_17 ), .B1(_10709_ ), .B2(_10710_ ), .ZN(_00429_ ) );
NAND4_X1 _14521_ ( .A1(_10263_ ), .A2(_10683_ ), .A3(_10684_ ), .A4(_09998_ ), .ZN(_10711_ ) );
OAI21_X1 _14522_ ( .A(\u_lsu.pmem[3878] ), .B1(_10257_ ), .B2(_10518_ ), .ZN(_10712_ ) );
AOI21_X1 _14523_ ( .A(fanout_net_17 ), .B1(_10711_ ), .B2(_10712_ ), .ZN(_00430_ ) );
OAI21_X1 _14524_ ( .A(\u_lsu.pmem[7552] ), .B1(_10692_ ), .B2(_10701_ ), .ZN(_10713_ ) );
NAND4_X1 _14525_ ( .A1(_10695_ ), .A2(_09548_ ), .A3(_10707_ ), .A4(_10461_ ), .ZN(_10714_ ) );
AOI21_X1 _14526_ ( .A(fanout_net_17 ), .B1(_10713_ ), .B2(_10714_ ), .ZN(_00431_ ) );
BUF_X4 _14527_ ( .A(_09108_ ), .Z(_10715_ ) );
NAND3_X1 _14528_ ( .A1(_10286_ ), .A2(_09558_ ), .A3(_09605_ ), .ZN(_10716_ ) );
NOR2_X1 _14529_ ( .A1(_09496_ ), .A2(_10716_ ), .ZN(_10717_ ) );
OAI21_X1 _14530_ ( .A(_10715_ ), .B1(_10717_ ), .B2(\u_lsu.pmem[7527] ), .ZN(_10718_ ) );
AOI21_X1 _14531_ ( .A(_10718_ ), .B1(_09638_ ), .B2(_10717_ ), .ZN(_00432_ ) );
BUF_X4 _14532_ ( .A(_09578_ ), .Z(_10719_ ) );
BUF_X4 _14533_ ( .A(_09450_ ), .Z(_10720_ ) );
BUF_X4 _14534_ ( .A(_10720_ ), .Z(_10721_ ) );
AND2_X1 _14535_ ( .A1(_10286_ ), .A2(_09558_ ), .ZN(_10722_ ) );
BUF_X4 _14536_ ( .A(_10722_ ), .Z(_10723_ ) );
BUF_X4 _14537_ ( .A(_10723_ ), .Z(_10724_ ) );
NAND4_X1 _14538_ ( .A1(_10719_ ), .A2(_10721_ ), .A3(_10684_ ), .A4(_10724_ ), .ZN(_10725_ ) );
BUF_X4 _14539_ ( .A(_10716_ ), .Z(_10726_ ) );
OAI21_X1 _14540_ ( .A(\u_lsu.pmem[7526] ), .B1(_10108_ ), .B2(_10726_ ), .ZN(_10727_ ) );
AOI21_X1 _14541_ ( .A(fanout_net_17 ), .B1(_10725_ ), .B2(_10727_ ), .ZN(_00433_ ) );
BUF_X4 _14542_ ( .A(_09585_ ), .Z(_10728_ ) );
NAND4_X1 _14543_ ( .A1(_10728_ ), .A2(_10721_ ), .A3(_10684_ ), .A4(_10724_ ), .ZN(_10729_ ) );
OAI21_X1 _14544_ ( .A(\u_lsu.pmem[7525] ), .B1(_10108_ ), .B2(_10726_ ), .ZN(_10730_ ) );
AOI21_X1 _14545_ ( .A(fanout_net_17 ), .B1(_10729_ ), .B2(_10730_ ), .ZN(_00434_ ) );
NAND4_X1 _14546_ ( .A1(_09589_ ), .A2(_10721_ ), .A3(_10684_ ), .A4(_10724_ ), .ZN(_10731_ ) );
OAI21_X1 _14547_ ( .A(\u_lsu.pmem[7524] ), .B1(_10108_ ), .B2(_10726_ ), .ZN(_10732_ ) );
AOI21_X1 _14548_ ( .A(fanout_net_17 ), .B1(_10731_ ), .B2(_10732_ ), .ZN(_00435_ ) );
BUF_X4 _14549_ ( .A(_09448_ ), .Z(_10733_ ) );
NAND4_X1 _14550_ ( .A1(_10733_ ), .A2(_10721_ ), .A3(_10684_ ), .A4(_10724_ ), .ZN(_10734_ ) );
OAI21_X1 _14551_ ( .A(\u_lsu.pmem[7523] ), .B1(_10108_ ), .B2(_10716_ ), .ZN(_10735_ ) );
AOI21_X1 _14552_ ( .A(fanout_net_17 ), .B1(_10734_ ), .B2(_10735_ ), .ZN(_00436_ ) );
NAND4_X1 _14553_ ( .A1(_09612_ ), .A2(_10721_ ), .A3(_10684_ ), .A4(_10724_ ), .ZN(_10736_ ) );
OAI21_X1 _14554_ ( .A(\u_lsu.pmem[7522] ), .B1(_10108_ ), .B2(_10716_ ), .ZN(_10737_ ) );
AOI21_X1 _14555_ ( .A(fanout_net_17 ), .B1(_10736_ ), .B2(_10737_ ), .ZN(_00437_ ) );
BUF_X4 _14556_ ( .A(_09616_ ), .Z(_10738_ ) );
NAND4_X1 _14557_ ( .A1(_10738_ ), .A2(_10721_ ), .A3(_10684_ ), .A4(_10724_ ), .ZN(_10739_ ) );
OAI21_X1 _14558_ ( .A(\u_lsu.pmem[7521] ), .B1(_10108_ ), .B2(_10716_ ), .ZN(_10740_ ) );
AOI21_X1 _14559_ ( .A(fanout_net_17 ), .B1(_10739_ ), .B2(_10740_ ), .ZN(_00438_ ) );
BUF_X4 _14560_ ( .A(_09621_ ), .Z(_10741_ ) );
NAND4_X1 _14561_ ( .A1(_10741_ ), .A2(_10721_ ), .A3(_10684_ ), .A4(_10724_ ), .ZN(_10742_ ) );
OAI21_X1 _14562_ ( .A(\u_lsu.pmem[7520] ), .B1(_10108_ ), .B2(_10716_ ), .ZN(_10743_ ) );
AOI21_X1 _14563_ ( .A(fanout_net_17 ), .B1(_10742_ ), .B2(_10743_ ), .ZN(_00439_ ) );
BUF_X2 _14564_ ( .A(_08993_ ), .Z(_10744_ ) );
AND2_X1 _14565_ ( .A1(_10744_ ), .A2(_09631_ ), .ZN(_10745_ ) );
AND2_X1 _14566_ ( .A1(_10745_ ), .A2(_09491_ ), .ZN(_10746_ ) );
INV_X1 _14567_ ( .A(_10746_ ), .ZN(_10747_ ) );
BUF_X4 _14568_ ( .A(_10747_ ), .Z(_10748_ ) );
OAI21_X1 _14569_ ( .A(\u_lsu.pmem[7495] ), .B1(_10748_ ), .B2(_10572_ ), .ZN(_10749_ ) );
BUF_X4 _14570_ ( .A(_10745_ ), .Z(_10750_ ) );
BUF_X4 _14571_ ( .A(_10750_ ), .Z(_10751_ ) );
BUF_X4 _14572_ ( .A(_08582_ ), .Z(_10752_ ) );
NAND4_X1 _14573_ ( .A1(_10751_ ), .A2(_10752_ ), .A3(_10589_ ), .A4(_10273_ ), .ZN(_10753_ ) );
AOI21_X1 _14574_ ( .A(fanout_net_17 ), .B1(_10749_ ), .B2(_10753_ ), .ZN(_00440_ ) );
NAND4_X1 _14575_ ( .A1(_10267_ ), .A2(_10683_ ), .A3(_10684_ ), .A4(_09998_ ), .ZN(_10754_ ) );
OAI21_X1 _14576_ ( .A(\u_lsu.pmem[3877] ), .B1(_10257_ ), .B2(_10518_ ), .ZN(_10755_ ) );
AOI21_X1 _14577_ ( .A(fanout_net_17 ), .B1(_10754_ ), .B2(_10755_ ), .ZN(_00441_ ) );
BUF_X4 _14578_ ( .A(_10340_ ), .Z(_10756_ ) );
NAND4_X1 _14579_ ( .A1(_10719_ ), .A2(_10721_ ), .A3(_10756_ ), .A4(_10751_ ), .ZN(_10757_ ) );
OAI21_X1 _14580_ ( .A(\u_lsu.pmem[7494] ), .B1(_10748_ ), .B2(_10140_ ), .ZN(_10758_ ) );
AOI21_X1 _14581_ ( .A(fanout_net_17 ), .B1(_10757_ ), .B2(_10758_ ), .ZN(_00442_ ) );
NAND4_X1 _14582_ ( .A1(_10728_ ), .A2(_10721_ ), .A3(_10756_ ), .A4(_10751_ ), .ZN(_10759_ ) );
BUF_X4 _14583_ ( .A(_10070_ ), .Z(_10760_ ) );
OAI21_X1 _14584_ ( .A(\u_lsu.pmem[7493] ), .B1(_10748_ ), .B2(_10760_ ), .ZN(_10761_ ) );
AOI21_X1 _14585_ ( .A(fanout_net_17 ), .B1(_10759_ ), .B2(_10761_ ), .ZN(_00443_ ) );
NAND4_X1 _14586_ ( .A1(_09589_ ), .A2(_10721_ ), .A3(_10756_ ), .A4(_10751_ ), .ZN(_10762_ ) );
OAI21_X1 _14587_ ( .A(\u_lsu.pmem[7492] ), .B1(_10748_ ), .B2(_10760_ ), .ZN(_10763_ ) );
AOI21_X1 _14588_ ( .A(fanout_net_17 ), .B1(_10762_ ), .B2(_10763_ ), .ZN(_00444_ ) );
NAND4_X1 _14589_ ( .A1(_10733_ ), .A2(_10034_ ), .A3(_10756_ ), .A4(_10751_ ), .ZN(_10764_ ) );
OAI21_X1 _14590_ ( .A(\u_lsu.pmem[7491] ), .B1(_10748_ ), .B2(_10760_ ), .ZN(_10765_ ) );
AOI21_X1 _14591_ ( .A(fanout_net_17 ), .B1(_10764_ ), .B2(_10765_ ), .ZN(_00445_ ) );
NAND4_X1 _14592_ ( .A1(_09612_ ), .A2(_10034_ ), .A3(_10756_ ), .A4(_10751_ ), .ZN(_10766_ ) );
OAI21_X1 _14593_ ( .A(\u_lsu.pmem[7490] ), .B1(_10748_ ), .B2(_10760_ ), .ZN(_10767_ ) );
AOI21_X1 _14594_ ( .A(fanout_net_17 ), .B1(_10766_ ), .B2(_10767_ ), .ZN(_00446_ ) );
NAND4_X1 _14595_ ( .A1(_10738_ ), .A2(_10034_ ), .A3(_10756_ ), .A4(_10751_ ), .ZN(_10768_ ) );
OAI21_X1 _14596_ ( .A(\u_lsu.pmem[7489] ), .B1(_10748_ ), .B2(_10760_ ), .ZN(_10769_ ) );
AOI21_X1 _14597_ ( .A(fanout_net_17 ), .B1(_10768_ ), .B2(_10769_ ), .ZN(_00447_ ) );
NAND4_X1 _14598_ ( .A1(_09622_ ), .A2(_10034_ ), .A3(_10756_ ), .A4(_10751_ ), .ZN(_10770_ ) );
OAI21_X1 _14599_ ( .A(\u_lsu.pmem[7488] ), .B1(_10748_ ), .B2(_10760_ ), .ZN(_10771_ ) );
AOI21_X1 _14600_ ( .A(fanout_net_17 ), .B1(_10770_ ), .B2(_10771_ ), .ZN(_00448_ ) );
NAND4_X1 _14601_ ( .A1(_09670_ ), .A2(_10683_ ), .A3(_10756_ ), .A4(_10685_ ), .ZN(_10772_ ) );
AND3_X2 _14602_ ( .A1(_09118_ ), .A2(_09127_ ), .A3(_09129_ ), .ZN(_10773_ ) );
AND2_X2 _14603_ ( .A1(_10773_ ), .A2(_10325_ ), .ZN(_10774_ ) );
INV_X1 _14604_ ( .A(_10774_ ), .ZN(_10775_ ) );
BUF_X4 _14605_ ( .A(_10775_ ), .Z(_10776_ ) );
OAI21_X1 _14606_ ( .A(\u_lsu.pmem[7463] ), .B1(_10776_ ), .B2(_10465_ ), .ZN(_10777_ ) );
AOI21_X1 _14607_ ( .A(fanout_net_17 ), .B1(_10772_ ), .B2(_10777_ ), .ZN(_00449_ ) );
NAND4_X1 _14608_ ( .A1(_09681_ ), .A2(_10683_ ), .A3(_10756_ ), .A4(_10685_ ), .ZN(_10778_ ) );
OAI21_X1 _14609_ ( .A(\u_lsu.pmem[7462] ), .B1(_10776_ ), .B2(_10465_ ), .ZN(_10779_ ) );
AOI21_X1 _14610_ ( .A(fanout_net_17 ), .B1(_10778_ ), .B2(_10779_ ), .ZN(_00450_ ) );
NAND4_X1 _14611_ ( .A1(_09685_ ), .A2(_10683_ ), .A3(_10756_ ), .A4(_10685_ ), .ZN(_10780_ ) );
OAI21_X1 _14612_ ( .A(\u_lsu.pmem[7461] ), .B1(_10775_ ), .B2(_10465_ ), .ZN(_10781_ ) );
AOI21_X1 _14613_ ( .A(fanout_net_17 ), .B1(_10780_ ), .B2(_10781_ ), .ZN(_00451_ ) );
AND2_X1 _14614_ ( .A1(_10255_ ), .A2(_10012_ ), .ZN(_10782_ ) );
OAI21_X1 _14615_ ( .A(_10715_ ), .B1(_10782_ ), .B2(\u_lsu.pmem[3876] ), .ZN(_10783_ ) );
AOI21_X1 _14616_ ( .A(_10783_ ), .B1(_09691_ ), .B2(_10782_ ), .ZN(_00452_ ) );
OAI21_X1 _14617_ ( .A(\u_lsu.pmem[7460] ), .B1(_10776_ ), .B2(_10701_ ), .ZN(_10784_ ) );
BUF_X4 _14618_ ( .A(_09472_ ), .Z(_10785_ ) );
NAND3_X1 _14619_ ( .A1(_10774_ ), .A2(_09589_ ), .A3(_10785_ ), .ZN(_10786_ ) );
AOI21_X1 _14620_ ( .A(fanout_net_17 ), .B1(_10784_ ), .B2(_10786_ ), .ZN(_00453_ ) );
OAI21_X1 _14621_ ( .A(\u_lsu.pmem[7459] ), .B1(_10776_ ), .B2(_10701_ ), .ZN(_10787_ ) );
NAND3_X1 _14622_ ( .A1(_10774_ ), .A2(_09592_ ), .A3(_10785_ ), .ZN(_10788_ ) );
AOI21_X1 _14623_ ( .A(fanout_net_17 ), .B1(_10787_ ), .B2(_10788_ ), .ZN(_00454_ ) );
OAI21_X1 _14624_ ( .A(\u_lsu.pmem[7458] ), .B1(_10776_ ), .B2(_10701_ ), .ZN(_10789_ ) );
NAND3_X1 _14625_ ( .A1(_10774_ ), .A2(_09695_ ), .A3(_10785_ ), .ZN(_10790_ ) );
AOI21_X1 _14626_ ( .A(fanout_net_17 ), .B1(_10789_ ), .B2(_10790_ ), .ZN(_00455_ ) );
OAI21_X1 _14627_ ( .A(\u_lsu.pmem[7457] ), .B1(_10776_ ), .B2(_10701_ ), .ZN(_10791_ ) );
NAND3_X1 _14628_ ( .A1(_10774_ ), .A2(_09617_ ), .A3(_10785_ ), .ZN(_10792_ ) );
AOI21_X1 _14629_ ( .A(fanout_net_17 ), .B1(_10791_ ), .B2(_10792_ ), .ZN(_00456_ ) );
BUF_X4 _14630_ ( .A(_10340_ ), .Z(_10793_ ) );
NAND4_X1 _14631_ ( .A1(_09703_ ), .A2(_10683_ ), .A3(_10793_ ), .A4(_10685_ ), .ZN(_10794_ ) );
OAI21_X1 _14632_ ( .A(\u_lsu.pmem[7456] ), .B1(_10775_ ), .B2(_10465_ ), .ZN(_10795_ ) );
AOI21_X1 _14633_ ( .A(fanout_net_18 ), .B1(_10794_ ), .B2(_10795_ ), .ZN(_00457_ ) );
NAND4_X1 _14634_ ( .A1(_09708_ ), .A2(_10636_ ), .A3(_10642_ ), .A4(_10646_ ), .ZN(_10796_ ) );
AND3_X1 _14635_ ( .A1(_09118_ ), .A2(_09505_ ), .A3(_09465_ ), .ZN(_10797_ ) );
NAND2_X4 _14636_ ( .A1(_10797_ ), .A2(_10326_ ), .ZN(_10798_ ) );
BUF_X4 _14637_ ( .A(_10798_ ), .Z(_10799_ ) );
OAI21_X1 _14638_ ( .A(\u_lsu.pmem[7431] ), .B1(_10660_ ), .B2(_10799_ ), .ZN(_10800_ ) );
AOI21_X1 _14639_ ( .A(fanout_net_18 ), .B1(_10796_ ), .B2(_10800_ ), .ZN(_00458_ ) );
NAND4_X1 _14640_ ( .A1(_09715_ ), .A2(_10636_ ), .A3(_10642_ ), .A4(_10646_ ), .ZN(_10801_ ) );
OAI21_X1 _14641_ ( .A(\u_lsu.pmem[7430] ), .B1(_10660_ ), .B2(_10799_ ), .ZN(_10802_ ) );
AOI21_X1 _14642_ ( .A(fanout_net_18 ), .B1(_10801_ ), .B2(_10802_ ), .ZN(_00459_ ) );
BUF_X4 _14643_ ( .A(_10585_ ), .Z(_10803_ ) );
NAND4_X1 _14644_ ( .A1(_09718_ ), .A2(_10803_ ), .A3(_10793_ ), .A4(_10685_ ), .ZN(_10804_ ) );
OAI21_X1 _14645_ ( .A(\u_lsu.pmem[7429] ), .B1(_10660_ ), .B2(_10799_ ), .ZN(_10805_ ) );
AOI21_X1 _14646_ ( .A(fanout_net_18 ), .B1(_10804_ ), .B2(_10805_ ), .ZN(_00460_ ) );
NAND4_X1 _14647_ ( .A1(_09721_ ), .A2(_10636_ ), .A3(_10642_ ), .A4(_10646_ ), .ZN(_10806_ ) );
BUF_X4 _14648_ ( .A(_10036_ ), .Z(_10807_ ) );
OAI21_X1 _14649_ ( .A(\u_lsu.pmem[7428] ), .B1(_10807_ ), .B2(_10799_ ), .ZN(_10808_ ) );
AOI21_X1 _14650_ ( .A(fanout_net_18 ), .B1(_10806_ ), .B2(_10808_ ), .ZN(_00461_ ) );
NAND4_X1 _14651_ ( .A1(_09725_ ), .A2(_10803_ ), .A3(_10793_ ), .A4(_10685_ ), .ZN(_10809_ ) );
OAI21_X1 _14652_ ( .A(\u_lsu.pmem[7427] ), .B1(_10807_ ), .B2(_10799_ ), .ZN(_10810_ ) );
AOI21_X1 _14653_ ( .A(fanout_net_18 ), .B1(_10809_ ), .B2(_10810_ ), .ZN(_00462_ ) );
OR4_X1 _14654_ ( .A1(_09969_ ), .A2(_10256_ ), .A3(_10045_ ), .A4(_10302_ ), .ZN(_10811_ ) );
OAI21_X1 _14655_ ( .A(\u_lsu.pmem[3875] ), .B1(_10256_ ), .B2(_10518_ ), .ZN(_10812_ ) );
AOI21_X1 _14656_ ( .A(fanout_net_18 ), .B1(_10811_ ), .B2(_10812_ ), .ZN(_00463_ ) );
OAI21_X1 _14657_ ( .A(\u_lsu.pmem[7426] ), .B1(_10546_ ), .B2(_10799_ ), .ZN(_10813_ ) );
NAND4_X1 _14658_ ( .A1(_09473_ ), .A2(_09474_ ), .A3(_10707_ ), .A4(_10797_ ), .ZN(_10814_ ) );
AOI21_X1 _14659_ ( .A(fanout_net_18 ), .B1(_10813_ ), .B2(_10814_ ), .ZN(_00464_ ) );
NAND4_X1 _14660_ ( .A1(_09733_ ), .A2(_10683_ ), .A3(_10793_ ), .A4(_10685_ ), .ZN(_10815_ ) );
OAI21_X1 _14661_ ( .A(\u_lsu.pmem[7425] ), .B1(_10807_ ), .B2(_10799_ ), .ZN(_10816_ ) );
AOI21_X1 _14662_ ( .A(fanout_net_18 ), .B1(_10815_ ), .B2(_10816_ ), .ZN(_00465_ ) );
NAND4_X1 _14663_ ( .A1(_09736_ ), .A2(_10636_ ), .A3(_10642_ ), .A4(_10646_ ), .ZN(_10817_ ) );
OAI21_X1 _14664_ ( .A(\u_lsu.pmem[7424] ), .B1(_10807_ ), .B2(_10799_ ), .ZN(_10818_ ) );
AOI21_X1 _14665_ ( .A(fanout_net_18 ), .B1(_10817_ ), .B2(_10818_ ), .ZN(_00466_ ) );
NOR2_X1 _14666_ ( .A1(_09506_ ), .A2(_09748_ ), .ZN(_10819_ ) );
NAND2_X1 _14667_ ( .A1(_10819_ ), .A2(_10326_ ), .ZN(_10820_ ) );
BUF_X4 _14668_ ( .A(_10820_ ), .Z(_10821_ ) );
OAI21_X1 _14669_ ( .A(\u_lsu.pmem[7399] ), .B1(_10546_ ), .B2(_10821_ ), .ZN(_10822_ ) );
NAND4_X1 _14670_ ( .A1(_10330_ ), .A2(_10549_ ), .A3(_10707_ ), .A4(_10819_ ), .ZN(_10823_ ) );
AOI21_X1 _14671_ ( .A(fanout_net_18 ), .B1(_10822_ ), .B2(_10823_ ), .ZN(_00467_ ) );
BUF_X4 _14672_ ( .A(_10046_ ), .Z(_10824_ ) );
NAND4_X1 _14673_ ( .A1(_09756_ ), .A2(_10824_ ), .A3(_10642_ ), .A4(_10646_ ), .ZN(_10825_ ) );
OAI21_X1 _14674_ ( .A(\u_lsu.pmem[7398] ), .B1(_10807_ ), .B2(_10821_ ), .ZN(_10826_ ) );
AOI21_X1 _14675_ ( .A(fanout_net_18 ), .B1(_10825_ ), .B2(_10826_ ), .ZN(_00468_ ) );
NAND4_X1 _14676_ ( .A1(_09763_ ), .A2(_10683_ ), .A3(_10793_ ), .A4(_10685_ ), .ZN(_10827_ ) );
OAI21_X1 _14677_ ( .A(\u_lsu.pmem[7397] ), .B1(_10807_ ), .B2(_10821_ ), .ZN(_10828_ ) );
AOI21_X1 _14678_ ( .A(fanout_net_18 ), .B1(_10827_ ), .B2(_10828_ ), .ZN(_00469_ ) );
NAND4_X1 _14679_ ( .A1(_09770_ ), .A2(_10803_ ), .A3(_10793_ ), .A4(_10685_ ), .ZN(_10829_ ) );
OAI21_X1 _14680_ ( .A(\u_lsu.pmem[7396] ), .B1(_10807_ ), .B2(_10821_ ), .ZN(_10830_ ) );
AOI21_X1 _14681_ ( .A(fanout_net_18 ), .B1(_10829_ ), .B2(_10830_ ), .ZN(_00470_ ) );
BUF_X4 _14682_ ( .A(_10592_ ), .Z(_10831_ ) );
NAND4_X1 _14683_ ( .A1(_09775_ ), .A2(_10683_ ), .A3(_10793_ ), .A4(_10831_ ), .ZN(_10832_ ) );
OAI21_X1 _14684_ ( .A(\u_lsu.pmem[7395] ), .B1(_10807_ ), .B2(_10821_ ), .ZN(_10833_ ) );
AOI21_X1 _14685_ ( .A(fanout_net_18 ), .B1(_10832_ ), .B2(_10833_ ), .ZN(_00471_ ) );
BUF_X4 _14686_ ( .A(_10126_ ), .Z(_10834_ ) );
NAND4_X1 _14687_ ( .A1(_09780_ ), .A2(_10834_ ), .A3(_10793_ ), .A4(_10831_ ), .ZN(_10835_ ) );
OAI21_X1 _14688_ ( .A(\u_lsu.pmem[7394] ), .B1(_10807_ ), .B2(_10821_ ), .ZN(_10836_ ) );
AOI21_X1 _14689_ ( .A(fanout_net_18 ), .B1(_10835_ ), .B2(_10836_ ), .ZN(_00472_ ) );
NAND4_X1 _14690_ ( .A1(_09787_ ), .A2(_10834_ ), .A3(_10793_ ), .A4(_10831_ ), .ZN(_10837_ ) );
OAI21_X1 _14691_ ( .A(\u_lsu.pmem[7393] ), .B1(_10807_ ), .B2(_10821_ ), .ZN(_10838_ ) );
AOI21_X1 _14692_ ( .A(fanout_net_18 ), .B1(_10837_ ), .B2(_10838_ ), .ZN(_00473_ ) );
OAI21_X1 _14693_ ( .A(\u_lsu.pmem[4327] ), .B1(_10546_ ), .B2(_09752_ ), .ZN(_10839_ ) );
NAND4_X1 _14694_ ( .A1(_10330_ ), .A2(_10549_ ), .A3(_09909_ ), .A4(_09749_ ), .ZN(_10840_ ) );
AOI21_X1 _14695_ ( .A(fanout_net_18 ), .B1(_10839_ ), .B2(_10840_ ), .ZN(_00474_ ) );
OR4_X1 _14696_ ( .A1(_09973_ ), .A2(_10256_ ), .A3(_10045_ ), .A4(_10302_ ), .ZN(_10841_ ) );
OAI21_X1 _14697_ ( .A(\u_lsu.pmem[3874] ), .B1(_10256_ ), .B2(_10518_ ), .ZN(_10842_ ) );
AOI21_X1 _14698_ ( .A(fanout_net_18 ), .B1(_10841_ ), .B2(_10842_ ), .ZN(_00475_ ) );
NAND4_X1 _14699_ ( .A1(_09791_ ), .A2(_10834_ ), .A3(_10793_ ), .A4(_10831_ ), .ZN(_10843_ ) );
BUF_X8 _14700_ ( .A(_09458_ ), .Z(_10844_ ) );
BUF_X4 _14701_ ( .A(_10844_ ), .Z(_10845_ ) );
OAI21_X1 _14702_ ( .A(\u_lsu.pmem[7392] ), .B1(_10845_ ), .B2(_10821_ ), .ZN(_10846_ ) );
AOI21_X1 _14703_ ( .A(fanout_net_18 ), .B1(_10843_ ), .B2(_10846_ ), .ZN(_00476_ ) );
NOR2_X1 _14704_ ( .A1(_09506_ ), .A2(_09797_ ), .ZN(_10847_ ) );
NAND2_X1 _14705_ ( .A1(_10847_ ), .A2(_10326_ ), .ZN(_10848_ ) );
BUF_X4 _14706_ ( .A(_10848_ ), .Z(_10849_ ) );
OAI21_X1 _14707_ ( .A(\u_lsu.pmem[7367] ), .B1(_10546_ ), .B2(_10849_ ), .ZN(_10850_ ) );
BUF_X4 _14708_ ( .A(_09741_ ), .Z(_10851_ ) );
NAND4_X1 _14709_ ( .A1(_10851_ ), .A2(_10549_ ), .A3(_10707_ ), .A4(_10847_ ), .ZN(_10852_ ) );
AOI21_X1 _14710_ ( .A(fanout_net_18 ), .B1(_10850_ ), .B2(_10852_ ), .ZN(_00477_ ) );
NAND4_X1 _14711_ ( .A1(_09804_ ), .A2(_10824_ ), .A3(\alu_result_out[8] ), .A4(_10585_ ), .ZN(_10853_ ) );
OAI21_X1 _14712_ ( .A(\u_lsu.pmem[7366] ), .B1(_10845_ ), .B2(_10849_ ), .ZN(_10854_ ) );
AOI21_X1 _14713_ ( .A(fanout_net_18 ), .B1(_10853_ ), .B2(_10854_ ), .ZN(_00478_ ) );
BUF_X4 _14714_ ( .A(_10340_ ), .Z(_10855_ ) );
NAND4_X1 _14715_ ( .A1(_09811_ ), .A2(_10803_ ), .A3(_10855_ ), .A4(_10831_ ), .ZN(_10856_ ) );
OAI21_X1 _14716_ ( .A(\u_lsu.pmem[7365] ), .B1(_10845_ ), .B2(_10849_ ), .ZN(_10857_ ) );
AOI21_X1 _14717_ ( .A(fanout_net_18 ), .B1(_10856_ ), .B2(_10857_ ), .ZN(_00479_ ) );
NAND4_X1 _14718_ ( .A1(_09815_ ), .A2(_10803_ ), .A3(_10855_ ), .A4(_10831_ ), .ZN(_10858_ ) );
OAI21_X1 _14719_ ( .A(\u_lsu.pmem[7364] ), .B1(_10845_ ), .B2(_10849_ ), .ZN(_10859_ ) );
AOI21_X1 _14720_ ( .A(fanout_net_18 ), .B1(_10858_ ), .B2(_10859_ ), .ZN(_00480_ ) );
NAND4_X1 _14721_ ( .A1(_09819_ ), .A2(_10803_ ), .A3(_10855_ ), .A4(_10831_ ), .ZN(_10860_ ) );
OAI21_X1 _14722_ ( .A(\u_lsu.pmem[7363] ), .B1(_10845_ ), .B2(_10849_ ), .ZN(_10861_ ) );
AOI21_X1 _14723_ ( .A(fanout_net_18 ), .B1(_10860_ ), .B2(_10861_ ), .ZN(_00481_ ) );
NAND4_X1 _14724_ ( .A1(_09827_ ), .A2(_10834_ ), .A3(_10855_ ), .A4(_10831_ ), .ZN(_10862_ ) );
OAI21_X1 _14725_ ( .A(\u_lsu.pmem[7362] ), .B1(_10845_ ), .B2(_10849_ ), .ZN(_10863_ ) );
AOI21_X1 _14726_ ( .A(fanout_net_18 ), .B1(_10862_ ), .B2(_10863_ ), .ZN(_00482_ ) );
NAND4_X1 _14727_ ( .A1(_09831_ ), .A2(_10834_ ), .A3(_10855_ ), .A4(_10831_ ), .ZN(_10864_ ) );
OAI21_X1 _14728_ ( .A(\u_lsu.pmem[7361] ), .B1(_10845_ ), .B2(_10849_ ), .ZN(_10865_ ) );
AOI21_X1 _14729_ ( .A(fanout_net_18 ), .B1(_10864_ ), .B2(_10865_ ), .ZN(_00483_ ) );
NAND4_X1 _14730_ ( .A1(_09835_ ), .A2(_10834_ ), .A3(_10855_ ), .A4(_10831_ ), .ZN(_10866_ ) );
OAI21_X1 _14731_ ( .A(\u_lsu.pmem[7360] ), .B1(_10845_ ), .B2(_10849_ ), .ZN(_10867_ ) );
AOI21_X1 _14732_ ( .A(fanout_net_18 ), .B1(_10866_ ), .B2(_10867_ ), .ZN(_00484_ ) );
BUF_X4 _14733_ ( .A(_10592_ ), .Z(_10868_ ) );
NAND4_X1 _14734_ ( .A1(_09840_ ), .A2(_10834_ ), .A3(_10855_ ), .A4(_10868_ ), .ZN(_10869_ ) );
NAND3_X1 _14735_ ( .A1(_10424_ ), .A2(_09743_ ), .A3(_09844_ ), .ZN(_10870_ ) );
BUF_X4 _14736_ ( .A(_10870_ ), .Z(_10871_ ) );
OAI21_X1 _14737_ ( .A(\u_lsu.pmem[7335] ), .B1(_10845_ ), .B2(_10871_ ), .ZN(_10872_ ) );
AOI21_X1 _14738_ ( .A(fanout_net_18 ), .B1(_10869_ ), .B2(_10872_ ), .ZN(_00485_ ) );
CLKBUF_X2 _14739_ ( .A(_09137_ ), .Z(_10873_ ) );
OR4_X1 _14740_ ( .A1(_09977_ ), .A2(_10256_ ), .A3(_10045_ ), .A4(_10873_ ), .ZN(_10874_ ) );
OAI21_X1 _14741_ ( .A(\u_lsu.pmem[3873] ), .B1(_10256_ ), .B2(_10518_ ), .ZN(_10875_ ) );
AOI21_X1 _14742_ ( .A(fanout_net_18 ), .B1(_10874_ ), .B2(_10875_ ), .ZN(_00486_ ) );
BUF_X4 _14743_ ( .A(_10287_ ), .Z(_10876_ ) );
NAND4_X1 _14744_ ( .A1(_09849_ ), .A2(_10824_ ), .A3(_10876_ ), .A4(_10646_ ), .ZN(_10877_ ) );
OAI21_X1 _14745_ ( .A(\u_lsu.pmem[7334] ), .B1(_10845_ ), .B2(_10871_ ), .ZN(_10878_ ) );
AOI21_X1 _14746_ ( .A(fanout_net_19 ), .B1(_10877_ ), .B2(_10878_ ), .ZN(_00487_ ) );
NAND4_X1 _14747_ ( .A1(_09853_ ), .A2(_10834_ ), .A3(_10855_ ), .A4(_10868_ ), .ZN(_10879_ ) );
BUF_X4 _14748_ ( .A(_10844_ ), .Z(_10880_ ) );
OAI21_X1 _14749_ ( .A(\u_lsu.pmem[7333] ), .B1(_10880_ ), .B2(_10871_ ), .ZN(_10881_ ) );
AOI21_X1 _14750_ ( .A(fanout_net_19 ), .B1(_10879_ ), .B2(_10881_ ), .ZN(_00488_ ) );
NAND4_X1 _14751_ ( .A1(_09858_ ), .A2(_10834_ ), .A3(_10855_ ), .A4(_10868_ ), .ZN(_10882_ ) );
OAI21_X1 _14752_ ( .A(\u_lsu.pmem[7332] ), .B1(_10880_ ), .B2(_10871_ ), .ZN(_10883_ ) );
AOI21_X1 _14753_ ( .A(fanout_net_19 ), .B1(_10882_ ), .B2(_10883_ ), .ZN(_00489_ ) );
NAND4_X1 _14754_ ( .A1(_09861_ ), .A2(_10834_ ), .A3(_10855_ ), .A4(_10868_ ), .ZN(_10884_ ) );
OAI21_X1 _14755_ ( .A(\u_lsu.pmem[7331] ), .B1(_10880_ ), .B2(_10871_ ), .ZN(_10885_ ) );
AOI21_X1 _14756_ ( .A(fanout_net_19 ), .B1(_10884_ ), .B2(_10885_ ), .ZN(_00490_ ) );
BUF_X8 _14757_ ( .A(_09875_ ), .Z(_10886_ ) );
BUF_X4 _14758_ ( .A(_10886_ ), .Z(_10887_ ) );
BUF_X4 _14759_ ( .A(_10340_ ), .Z(_10888_ ) );
NAND4_X1 _14760_ ( .A1(_09864_ ), .A2(_10887_ ), .A3(_10888_ ), .A4(_10868_ ), .ZN(_10889_ ) );
OAI21_X1 _14761_ ( .A(\u_lsu.pmem[7330] ), .B1(_10880_ ), .B2(_10871_ ), .ZN(_10890_ ) );
AOI21_X1 _14762_ ( .A(fanout_net_19 ), .B1(_10889_ ), .B2(_10890_ ), .ZN(_00491_ ) );
NAND4_X1 _14763_ ( .A1(_09867_ ), .A2(_10887_ ), .A3(_10888_ ), .A4(_10868_ ), .ZN(_10891_ ) );
OAI21_X1 _14764_ ( .A(\u_lsu.pmem[7329] ), .B1(_10880_ ), .B2(_10871_ ), .ZN(_10892_ ) );
AOI21_X1 _14765_ ( .A(fanout_net_19 ), .B1(_10891_ ), .B2(_10892_ ), .ZN(_00492_ ) );
NAND4_X1 _14766_ ( .A1(_09881_ ), .A2(_10803_ ), .A3(_10888_ ), .A4(_10868_ ), .ZN(_10893_ ) );
OAI21_X1 _14767_ ( .A(\u_lsu.pmem[7328] ), .B1(_10880_ ), .B2(_10871_ ), .ZN(_10894_ ) );
AOI21_X1 _14768_ ( .A(fanout_net_19 ), .B1(_10893_ ), .B2(_10894_ ), .ZN(_00493_ ) );
OR3_X4 _14769_ ( .A1(_09889_ ), .A2(_09842_ ), .A3(_09454_ ), .ZN(_10895_ ) );
BUF_X4 _14770_ ( .A(_10895_ ), .Z(_10896_ ) );
OAI21_X1 _14771_ ( .A(\u_lsu.pmem[7303] ), .B1(_10896_ ), .B2(_10701_ ), .ZN(_10897_ ) );
NOR2_X2 _14772_ ( .A1(_09889_ ), .A2(_09539_ ), .ZN(_10898_ ) );
BUF_X4 _14773_ ( .A(_10898_ ), .Z(_10899_ ) );
NAND4_X1 _14774_ ( .A1(_10899_ ), .A2(_10752_ ), .A3(_10707_ ), .A4(_10461_ ), .ZN(_10900_ ) );
AOI21_X1 _14775_ ( .A(fanout_net_19 ), .B1(_10897_ ), .B2(_10900_ ), .ZN(_00494_ ) );
BUF_X8 _14776_ ( .A(_09442_ ), .Z(_10901_ ) );
BUF_X4 _14777_ ( .A(_10901_ ), .Z(_10902_ ) );
OAI21_X1 _14778_ ( .A(\u_lsu.pmem[7302] ), .B1(_10896_ ), .B2(_10902_ ), .ZN(_10903_ ) );
BUF_X8 _14779_ ( .A(_09450_ ), .Z(_10904_ ) );
BUF_X4 _14780_ ( .A(_10904_ ), .Z(_10905_ ) );
NAND4_X1 _14781_ ( .A1(_10899_ ), .A2(_10185_ ), .A3(_10707_ ), .A4(_10905_ ), .ZN(_10906_ ) );
AOI21_X1 _14782_ ( .A(fanout_net_19 ), .B1(_10903_ ), .B2(_10906_ ), .ZN(_00495_ ) );
OAI21_X1 _14783_ ( .A(\u_lsu.pmem[7301] ), .B1(_10896_ ), .B2(_10902_ ), .ZN(_10907_ ) );
NAND4_X1 _14784_ ( .A1(_10899_ ), .A2(_10188_ ), .A3(_10707_ ), .A4(_10905_ ), .ZN(_10908_ ) );
AOI21_X1 _14785_ ( .A(fanout_net_19 ), .B1(_10907_ ), .B2(_10908_ ), .ZN(_00496_ ) );
NAND4_X1 _14786_ ( .A1(_10279_ ), .A2(_10887_ ), .A3(_10888_ ), .A4(_09998_ ), .ZN(_10909_ ) );
BUF_X4 _14787_ ( .A(_10046_ ), .Z(_10910_ ) );
OAI21_X1 _14788_ ( .A(\u_lsu.pmem[3872] ), .B1(_10256_ ), .B2(_10910_ ), .ZN(_10911_ ) );
AOI21_X1 _14789_ ( .A(fanout_net_19 ), .B1(_10909_ ), .B2(_10911_ ), .ZN(_00497_ ) );
OAI21_X1 _14790_ ( .A(\u_lsu.pmem[7300] ), .B1(_10896_ ), .B2(_10902_ ), .ZN(_10912_ ) );
NAND4_X1 _14791_ ( .A1(_10899_ ), .A2(_10192_ ), .A3(_10707_ ), .A4(_10905_ ), .ZN(_10913_ ) );
AOI21_X1 _14792_ ( .A(fanout_net_19 ), .B1(_10912_ ), .B2(_10913_ ), .ZN(_00498_ ) );
OAI21_X1 _14793_ ( .A(\u_lsu.pmem[7299] ), .B1(_10896_ ), .B2(_10902_ ), .ZN(_10914_ ) );
BUF_X4 _14794_ ( .A(_08650_ ), .Z(_10915_ ) );
BUF_X4 _14795_ ( .A(_09878_ ), .Z(_10916_ ) );
NAND4_X1 _14796_ ( .A1(_10899_ ), .A2(_10915_ ), .A3(_10916_ ), .A4(_10905_ ), .ZN(_10917_ ) );
AOI21_X1 _14797_ ( .A(fanout_net_19 ), .B1(_10914_ ), .B2(_10917_ ), .ZN(_00499_ ) );
OAI21_X1 _14798_ ( .A(\u_lsu.pmem[7298] ), .B1(_10896_ ), .B2(_10902_ ), .ZN(_10918_ ) );
NAND4_X1 _14799_ ( .A1(_09906_ ), .A2(_10437_ ), .A3(_10916_ ), .A4(_10905_ ), .ZN(_10919_ ) );
AOI21_X1 _14800_ ( .A(fanout_net_19 ), .B1(_10918_ ), .B2(_10919_ ), .ZN(_00500_ ) );
OAI21_X1 _14801_ ( .A(\u_lsu.pmem[7297] ), .B1(_10896_ ), .B2(_10902_ ), .ZN(_10920_ ) );
NAND4_X1 _14802_ ( .A1(_10899_ ), .A2(_09923_ ), .A3(_10916_ ), .A4(_10905_ ), .ZN(_10921_ ) );
AOI21_X1 _14803_ ( .A(fanout_net_19 ), .B1(_10920_ ), .B2(_10921_ ), .ZN(_00501_ ) );
OAI21_X1 _14804_ ( .A(\u_lsu.pmem[7296] ), .B1(_10896_ ), .B2(_10902_ ), .ZN(_10922_ ) );
NAND4_X1 _14805_ ( .A1(_10899_ ), .A2(_09548_ ), .A3(_10916_ ), .A4(_10905_ ), .ZN(_10923_ ) );
AOI21_X1 _14806_ ( .A(fanout_net_19 ), .B1(_10922_ ), .B2(_10923_ ), .ZN(_00502_ ) );
AND2_X1 _14807_ ( .A1(_09915_ ), .A2(_10744_ ), .ZN(_10924_ ) );
AND2_X1 _14808_ ( .A1(_10924_ ), .A2(_09605_ ), .ZN(_10925_ ) );
INV_X1 _14809_ ( .A(_10925_ ), .ZN(_10926_ ) );
BUF_X4 _14810_ ( .A(_10926_ ), .Z(_10927_ ) );
OAI21_X1 _14811_ ( .A(\u_lsu.pmem[7271] ), .B1(_10927_ ), .B2(_10902_ ), .ZN(_10928_ ) );
BUF_X4 _14812_ ( .A(_10924_ ), .Z(_10929_ ) );
BUF_X4 _14813_ ( .A(_10929_ ), .Z(_10930_ ) );
NAND4_X1 _14814_ ( .A1(_10930_ ), .A2(_10752_ ), .A3(_10589_ ), .A4(_10273_ ), .ZN(_10931_ ) );
AOI21_X1 _14815_ ( .A(fanout_net_19 ), .B1(_10928_ ), .B2(_10931_ ), .ZN(_00503_ ) );
OAI21_X1 _14816_ ( .A(\u_lsu.pmem[7270] ), .B1(_10927_ ), .B2(_10902_ ), .ZN(_10932_ ) );
NAND4_X1 _14817_ ( .A1(_09579_ ), .A2(_10549_ ), .A3(_10916_ ), .A4(_10930_ ), .ZN(_10933_ ) );
AOI21_X1 _14818_ ( .A(fanout_net_19 ), .B1(_10932_ ), .B2(_10933_ ), .ZN(_00504_ ) );
OAI21_X1 _14819_ ( .A(\u_lsu.pmem[7269] ), .B1(_10927_ ), .B2(_10902_ ), .ZN(_10934_ ) );
NAND4_X1 _14820_ ( .A1(_09586_ ), .A2(_10549_ ), .A3(_10916_ ), .A4(_10930_ ), .ZN(_10935_ ) );
AOI21_X1 _14821_ ( .A(fanout_net_19 ), .B1(_10934_ ), .B2(_10935_ ), .ZN(_00505_ ) );
BUF_X4 _14822_ ( .A(_10901_ ), .Z(_10936_ ) );
OAI21_X1 _14823_ ( .A(\u_lsu.pmem[7268] ), .B1(_10927_ ), .B2(_10936_ ), .ZN(_10937_ ) );
BUF_X4 _14824_ ( .A(_10548_ ), .Z(_10938_ ) );
BUF_X4 _14825_ ( .A(_10924_ ), .Z(_10939_ ) );
NAND4_X1 _14826_ ( .A1(_10486_ ), .A2(_10938_ ), .A3(_10916_ ), .A4(_10939_ ), .ZN(_10940_ ) );
AOI21_X1 _14827_ ( .A(fanout_net_19 ), .B1(_10937_ ), .B2(_10940_ ), .ZN(_00506_ ) );
OAI21_X1 _14828_ ( .A(\u_lsu.pmem[7267] ), .B1(_10927_ ), .B2(_10936_ ), .ZN(_10941_ ) );
NAND4_X1 _14829_ ( .A1(_09449_ ), .A2(_10938_ ), .A3(_10916_ ), .A4(_10939_ ), .ZN(_10942_ ) );
AOI21_X1 _14830_ ( .A(fanout_net_19 ), .B1(_10941_ ), .B2(_10942_ ), .ZN(_00507_ ) );
NAND4_X1 _14831_ ( .A1(_10285_ ), .A2(_10803_ ), .A3(_10888_ ), .A4(_09998_ ), .ZN(_10943_ ) );
NAND2_X1 _14832_ ( .A1(_10291_ ), .A2(_10012_ ), .ZN(_10944_ ) );
NAND2_X1 _14833_ ( .A1(_10944_ ), .A2(\u_lsu.pmem[3847] ), .ZN(_10945_ ) );
AOI21_X1 _14834_ ( .A(fanout_net_19 ), .B1(_10943_ ), .B2(_10945_ ), .ZN(_00508_ ) );
OAI21_X1 _14835_ ( .A(\u_lsu.pmem[7266] ), .B1(_10927_ ), .B2(_10936_ ), .ZN(_10946_ ) );
NAND4_X1 _14836_ ( .A1(_10492_ ), .A2(_10938_ ), .A3(_10916_ ), .A4(_10939_ ), .ZN(_10947_ ) );
AOI21_X1 _14837_ ( .A(fanout_net_19 ), .B1(_10946_ ), .B2(_10947_ ), .ZN(_00509_ ) );
OAI21_X1 _14838_ ( .A(\u_lsu.pmem[7265] ), .B1(_10927_ ), .B2(_10936_ ), .ZN(_10948_ ) );
NAND4_X1 _14839_ ( .A1(_09698_ ), .A2(_10938_ ), .A3(_10916_ ), .A4(_10939_ ), .ZN(_10949_ ) );
AOI21_X1 _14840_ ( .A(fanout_net_19 ), .B1(_10948_ ), .B2(_10949_ ), .ZN(_00510_ ) );
OAI21_X1 _14841_ ( .A(\u_lsu.pmem[7264] ), .B1(_10927_ ), .B2(_10936_ ), .ZN(_10950_ ) );
BUF_X4 _14842_ ( .A(_09878_ ), .Z(_10951_ ) );
NAND4_X1 _14843_ ( .A1(_10525_ ), .A2(_10938_ ), .A3(_10951_ ), .A4(_10939_ ), .ZN(_10952_ ) );
AOI21_X1 _14844_ ( .A(fanout_net_19 ), .B1(_10950_ ), .B2(_10952_ ), .ZN(_00511_ ) );
AND2_X1 _14845_ ( .A1(_09948_ ), .A2(_09489_ ), .ZN(_10953_ ) );
AND2_X1 _14846_ ( .A1(_10953_ ), .A2(_09491_ ), .ZN(_10954_ ) );
INV_X1 _14847_ ( .A(_10954_ ), .ZN(_10955_ ) );
BUF_X4 _14848_ ( .A(_10955_ ), .Z(_10956_ ) );
OAI21_X1 _14849_ ( .A(\u_lsu.pmem[7239] ), .B1(_10956_ ), .B2(_10572_ ), .ZN(_10957_ ) );
NAND4_X1 _14850_ ( .A1(_10953_ ), .A2(_10752_ ), .A3(_10589_ ), .A4(_09606_ ), .ZN(_10958_ ) );
AOI21_X1 _14851_ ( .A(fanout_net_19 ), .B1(_10957_ ), .B2(_10958_ ), .ZN(_00512_ ) );
OAI21_X1 _14852_ ( .A(\u_lsu.pmem[7238] ), .B1(_10956_ ), .B2(_10572_ ), .ZN(_10959_ ) );
NAND4_X1 _14853_ ( .A1(_09957_ ), .A2(_10437_ ), .A3(_10951_ ), .A4(_10905_ ), .ZN(_10960_ ) );
AOI21_X1 _14854_ ( .A(fanout_net_19 ), .B1(_10959_ ), .B2(_10960_ ), .ZN(_00513_ ) );
OAI21_X1 _14855_ ( .A(\u_lsu.pmem[7237] ), .B1(_10956_ ), .B2(_10572_ ), .ZN(_10961_ ) );
NAND4_X1 _14856_ ( .A1(_09961_ ), .A2(_10437_ ), .A3(_10951_ ), .A4(_10905_ ), .ZN(_10962_ ) );
AOI21_X1 _14857_ ( .A(fanout_net_19 ), .B1(_10961_ ), .B2(_10962_ ), .ZN(_00514_ ) );
OAI21_X1 _14858_ ( .A(\u_lsu.pmem[7236] ), .B1(_10956_ ), .B2(_10572_ ), .ZN(_10963_ ) );
NAND4_X1 _14859_ ( .A1(_09966_ ), .A2(_10437_ ), .A3(_10951_ ), .A4(_10905_ ), .ZN(_10964_ ) );
AOI21_X1 _14860_ ( .A(fanout_net_19 ), .B1(_10963_ ), .B2(_10964_ ), .ZN(_00515_ ) );
OAI21_X1 _14861_ ( .A(\u_lsu.pmem[7235] ), .B1(_10956_ ), .B2(_10572_ ), .ZN(_10965_ ) );
BUF_X4 _14862_ ( .A(_10904_ ), .Z(_10966_ ) );
NAND4_X1 _14863_ ( .A1(_09970_ ), .A2(_10437_ ), .A3(_10951_ ), .A4(_10966_ ), .ZN(_10967_ ) );
AOI21_X1 _14864_ ( .A(fanout_net_19 ), .B1(_10965_ ), .B2(_10967_ ), .ZN(_00516_ ) );
OAI21_X1 _14865_ ( .A(\u_lsu.pmem[7234] ), .B1(_10956_ ), .B2(_10572_ ), .ZN(_10968_ ) );
NAND4_X1 _14866_ ( .A1(_09974_ ), .A2(_10437_ ), .A3(_10951_ ), .A4(_10966_ ), .ZN(_10969_ ) );
AOI21_X1 _14867_ ( .A(fanout_net_20 ), .B1(_10968_ ), .B2(_10969_ ), .ZN(_00517_ ) );
OAI21_X1 _14868_ ( .A(\u_lsu.pmem[7233] ), .B1(_10956_ ), .B2(_10572_ ), .ZN(_10970_ ) );
NAND4_X1 _14869_ ( .A1(_09978_ ), .A2(_10437_ ), .A3(_10951_ ), .A4(_10966_ ), .ZN(_10971_ ) );
AOI21_X1 _14870_ ( .A(fanout_net_20 ), .B1(_10970_ ), .B2(_10971_ ), .ZN(_00518_ ) );
NAND4_X1 _14871_ ( .A1(_10295_ ), .A2(_10803_ ), .A3(_10888_ ), .A4(_09998_ ), .ZN(_10972_ ) );
NAND2_X1 _14872_ ( .A1(_10944_ ), .A2(\u_lsu.pmem[3846] ), .ZN(_10973_ ) );
AOI21_X1 _14873_ ( .A(fanout_net_20 ), .B1(_10972_ ), .B2(_10973_ ), .ZN(_00519_ ) );
BUF_X4 _14874_ ( .A(_10070_ ), .Z(_10974_ ) );
OAI21_X1 _14875_ ( .A(\u_lsu.pmem[7232] ), .B1(_10956_ ), .B2(_10974_ ), .ZN(_10975_ ) );
BUF_X4 _14876_ ( .A(_10063_ ), .Z(_10976_ ) );
NAND4_X1 _14877_ ( .A1(_09982_ ), .A2(_10976_ ), .A3(_10951_ ), .A4(_10966_ ), .ZN(_10977_ ) );
AOI21_X1 _14878_ ( .A(fanout_net_20 ), .B1(_10975_ ), .B2(_10977_ ), .ZN(_00520_ ) );
NAND4_X1 _14879_ ( .A1(_09987_ ), .A2(_10887_ ), .A3(_10888_ ), .A4(_10868_ ), .ZN(_10978_ ) );
AND2_X2 _14880_ ( .A1(_09989_ ), .A2(_10055_ ), .ZN(_10979_ ) );
AND2_X1 _14881_ ( .A1(_10979_ ), .A2(_09605_ ), .ZN(_10980_ ) );
NAND2_X1 _14882_ ( .A1(_10980_ ), .A2(_09950_ ), .ZN(_10981_ ) );
NAND2_X1 _14883_ ( .A1(_10981_ ), .A2(\u_lsu.pmem[7207] ), .ZN(_10982_ ) );
AOI21_X1 _14884_ ( .A(fanout_net_20 ), .B1(_10978_ ), .B2(_10982_ ), .ZN(_00521_ ) );
NAND4_X1 _14885_ ( .A1(_09994_ ), .A2(_10887_ ), .A3(_10888_ ), .A4(_10868_ ), .ZN(_10983_ ) );
NAND2_X1 _14886_ ( .A1(_10981_ ), .A2(\u_lsu.pmem[7206] ), .ZN(_10984_ ) );
AOI21_X1 _14887_ ( .A(fanout_net_20 ), .B1(_10983_ ), .B2(_10984_ ), .ZN(_00522_ ) );
NAND4_X1 _14888_ ( .A1(_09997_ ), .A2(_10887_ ), .A3(_10888_ ), .A4(_10868_ ), .ZN(_10985_ ) );
NAND2_X1 _14889_ ( .A1(_10981_ ), .A2(\u_lsu.pmem[7205] ), .ZN(_10986_ ) );
AOI21_X1 _14890_ ( .A(fanout_net_20 ), .B1(_10985_ ), .B2(_10986_ ), .ZN(_00523_ ) );
NAND2_X1 _14891_ ( .A1(_10981_ ), .A2(\u_lsu.pmem[7204] ), .ZN(_10987_ ) );
BUF_X4 _14892_ ( .A(_10979_ ), .Z(_10988_ ) );
NAND4_X1 _14893_ ( .A1(_10486_ ), .A2(_10938_ ), .A3(_10951_ ), .A4(_10988_ ), .ZN(_10989_ ) );
AOI21_X1 _14894_ ( .A(fanout_net_20 ), .B1(_10987_ ), .B2(_10989_ ), .ZN(_00524_ ) );
NAND2_X1 _14895_ ( .A1(_10981_ ), .A2(\u_lsu.pmem[7203] ), .ZN(_10990_ ) );
NAND4_X1 _14896_ ( .A1(_09449_ ), .A2(_10938_ ), .A3(_10951_ ), .A4(_10988_ ), .ZN(_10991_ ) );
AOI21_X1 _14897_ ( .A(fanout_net_20 ), .B1(_10990_ ), .B2(_10991_ ), .ZN(_00525_ ) );
NAND2_X1 _14898_ ( .A1(_10981_ ), .A2(\u_lsu.pmem[7202] ), .ZN(_10992_ ) );
BUF_X4 _14899_ ( .A(_09878_ ), .Z(_10993_ ) );
NAND4_X1 _14900_ ( .A1(_10492_ ), .A2(_10938_ ), .A3(_10993_ ), .A4(_10988_ ), .ZN(_10994_ ) );
AOI21_X1 _14901_ ( .A(fanout_net_20 ), .B1(_10992_ ), .B2(_10994_ ), .ZN(_00526_ ) );
NAND2_X1 _14902_ ( .A1(_10981_ ), .A2(\u_lsu.pmem[7201] ), .ZN(_10995_ ) );
NAND4_X1 _14903_ ( .A1(_09698_ ), .A2(_10938_ ), .A3(_10993_ ), .A4(_10988_ ), .ZN(_10996_ ) );
AOI21_X1 _14904_ ( .A(fanout_net_20 ), .B1(_10995_ ), .B2(_10996_ ), .ZN(_00527_ ) );
BUF_X4 _14905_ ( .A(_10592_ ), .Z(_10997_ ) );
NAND4_X1 _14906_ ( .A1(_10021_ ), .A2(_10887_ ), .A3(_10888_ ), .A4(_10997_ ), .ZN(_10998_ ) );
NAND2_X1 _14907_ ( .A1(_10981_ ), .A2(\u_lsu.pmem[7200] ), .ZN(_10999_ ) );
AOI21_X1 _14908_ ( .A(fanout_net_20 ), .B1(_10998_ ), .B2(_10999_ ), .ZN(_00528_ ) );
BUF_X4 _14909_ ( .A(_09741_ ), .Z(_11000_ ) );
AND2_X1 _14910_ ( .A1(_09116_ ), .A2(_08993_ ), .ZN(_11001_ ) );
NAND4_X1 _14911_ ( .A1(_11000_ ), .A2(_10824_ ), .A3(\alu_result_out[8] ), .A4(_11001_ ), .ZN(_11002_ ) );
AND2_X2 _14912_ ( .A1(_11001_ ), .A2(_09018_ ), .ZN(_11003_ ) );
INV_X1 _14913_ ( .A(_11003_ ), .ZN(_11004_ ) );
BUF_X4 _14914_ ( .A(_11004_ ), .Z(_11005_ ) );
BUF_X4 _14915_ ( .A(_11005_ ), .Z(_11006_ ) );
OAI21_X1 _14916_ ( .A(\u_lsu.pmem[7175] ), .B1(_11006_ ), .B2(_10760_ ), .ZN(_11007_ ) );
AOI21_X1 _14917_ ( .A(fanout_net_20 ), .B1(_11002_ ), .B2(_11007_ ), .ZN(_00529_ ) );
BUF_X4 _14918_ ( .A(_10340_ ), .Z(_11008_ ) );
NAND4_X1 _14919_ ( .A1(_10299_ ), .A2(_10803_ ), .A3(_11008_ ), .A4(_09998_ ), .ZN(_11009_ ) );
NAND2_X1 _14920_ ( .A1(_10944_ ), .A2(\u_lsu.pmem[3845] ), .ZN(_11010_ ) );
AOI21_X1 _14921_ ( .A(fanout_net_20 ), .B1(_11009_ ), .B2(_11010_ ), .ZN(_00530_ ) );
CLKBUF_X2 _14922_ ( .A(_09493_ ), .Z(_11011_ ) );
OR4_X1 _14923_ ( .A1(_09576_ ), .A2(_11005_ ), .A3(_11011_ ), .A4(_10873_ ), .ZN(_11012_ ) );
OAI21_X1 _14924_ ( .A(\u_lsu.pmem[7174] ), .B1(_11006_ ), .B2(_10760_ ), .ZN(_11013_ ) );
AOI21_X1 _14925_ ( .A(fanout_net_20 ), .B1(_11012_ ), .B2(_11013_ ), .ZN(_00531_ ) );
OR4_X1 _14926_ ( .A1(_09583_ ), .A2(_11005_ ), .A3(_11011_ ), .A4(_10873_ ), .ZN(_11014_ ) );
OAI21_X1 _14927_ ( .A(\u_lsu.pmem[7173] ), .B1(_11006_ ), .B2(_10760_ ), .ZN(_11015_ ) );
AOI21_X1 _14928_ ( .A(fanout_net_20 ), .B1(_11014_ ), .B2(_11015_ ), .ZN(_00532_ ) );
OR4_X1 _14929_ ( .A1(_09146_ ), .A2(_11005_ ), .A3(_11011_ ), .A4(_10873_ ), .ZN(_11016_ ) );
OAI21_X1 _14930_ ( .A(\u_lsu.pmem[7172] ), .B1(_11006_ ), .B2(_10760_ ), .ZN(_11017_ ) );
AOI21_X1 _14931_ ( .A(fanout_net_20 ), .B1(_11016_ ), .B2(_11017_ ), .ZN(_00533_ ) );
OR4_X1 _14932_ ( .A1(_09969_ ), .A2(_11004_ ), .A3(_11011_ ), .A4(_10873_ ), .ZN(_11018_ ) );
BUF_X4 _14933_ ( .A(_10070_ ), .Z(_11019_ ) );
OAI21_X1 _14934_ ( .A(\u_lsu.pmem[7171] ), .B1(_11006_ ), .B2(_11019_ ), .ZN(_11020_ ) );
AOI21_X1 _14935_ ( .A(fanout_net_20 ), .B1(_11018_ ), .B2(_11020_ ), .ZN(_00534_ ) );
NOR2_X1 _14936_ ( .A1(_10583_ ), .A2(_10061_ ), .ZN(_11021_ ) );
NAND4_X1 _14937_ ( .A1(_11021_ ), .A2(_09868_ ), .A3(_11008_ ), .A4(_10997_ ), .ZN(_11022_ ) );
OAI21_X1 _14938_ ( .A(\u_lsu.pmem[7170] ), .B1(_11006_ ), .B2(_11019_ ), .ZN(_11023_ ) );
AOI21_X1 _14939_ ( .A(fanout_net_20 ), .B1(_11022_ ), .B2(_11023_ ), .ZN(_00535_ ) );
OR4_X1 _14940_ ( .A1(_09977_ ), .A2(_11004_ ), .A3(_11011_ ), .A4(_10873_ ), .ZN(_11024_ ) );
OAI21_X1 _14941_ ( .A(\u_lsu.pmem[7169] ), .B1(_11006_ ), .B2(_11019_ ), .ZN(_11025_ ) );
AOI21_X1 _14942_ ( .A(fanout_net_20 ), .B1(_11024_ ), .B2(_11025_ ), .ZN(_00536_ ) );
OR4_X1 _14943_ ( .A1(_09497_ ), .A2(_11004_ ), .A3(_11011_ ), .A4(_10873_ ), .ZN(_11026_ ) );
OAI21_X1 _14944_ ( .A(\u_lsu.pmem[7168] ), .B1(_11006_ ), .B2(_11019_ ), .ZN(_11027_ ) );
AOI21_X1 _14945_ ( .A(fanout_net_20 ), .B1(_11026_ ), .B2(_11027_ ), .ZN(_00537_ ) );
BUF_X4 _14946_ ( .A(_10325_ ), .Z(_11028_ ) );
INV_X1 _14947_ ( .A(_10052_ ), .ZN(_11029_ ) );
NOR3_X4 _14948_ ( .A1(_10055_ ), .A2(_11029_ ), .A3(_09666_ ), .ZN(_11030_ ) );
NAND2_X1 _14949_ ( .A1(_11028_ ), .A2(_11030_ ), .ZN(_11031_ ) );
BUF_X4 _14950_ ( .A(_11031_ ), .Z(_11032_ ) );
OAI21_X1 _14951_ ( .A(\u_lsu.pmem[7143] ), .B1(_10546_ ), .B2(_11032_ ), .ZN(_11033_ ) );
NAND4_X1 _14952_ ( .A1(_10851_ ), .A2(_10938_ ), .A3(_10993_ ), .A4(_11030_ ), .ZN(_11034_ ) );
AOI21_X1 _14953_ ( .A(fanout_net_20 ), .B1(_11033_ ), .B2(_11034_ ), .ZN(_00538_ ) );
NAND4_X1 _14954_ ( .A1(_10062_ ), .A2(_09868_ ), .A3(_11008_ ), .A4(_10997_ ), .ZN(_11035_ ) );
OAI21_X1 _14955_ ( .A(\u_lsu.pmem[7142] ), .B1(_10880_ ), .B2(_11032_ ), .ZN(_11036_ ) );
AOI21_X1 _14956_ ( .A(fanout_net_20 ), .B1(_11035_ ), .B2(_11036_ ), .ZN(_00539_ ) );
NAND4_X1 _14957_ ( .A1(_10075_ ), .A2(_09868_ ), .A3(_11008_ ), .A4(_10997_ ), .ZN(_11037_ ) );
OAI21_X1 _14958_ ( .A(\u_lsu.pmem[7141] ), .B1(_10880_ ), .B2(_11032_ ), .ZN(_11038_ ) );
AOI21_X1 _14959_ ( .A(fanout_net_20 ), .B1(_11037_ ), .B2(_11038_ ), .ZN(_00540_ ) );
BUF_X4 _14960_ ( .A(_10585_ ), .Z(_11039_ ) );
NAND4_X1 _14961_ ( .A1(_10306_ ), .A2(_11039_ ), .A3(_11008_ ), .A4(_09998_ ), .ZN(_11040_ ) );
NAND2_X1 _14962_ ( .A1(_10944_ ), .A2(\u_lsu.pmem[3844] ), .ZN(_11041_ ) );
AOI21_X1 _14963_ ( .A(fanout_net_20 ), .B1(_11040_ ), .B2(_11041_ ), .ZN(_00541_ ) );
BUF_X4 _14964_ ( .A(_09671_ ), .Z(_11042_ ) );
NAND4_X1 _14965_ ( .A1(_10079_ ), .A2(_11042_ ), .A3(_11008_ ), .A4(_10997_ ), .ZN(_11043_ ) );
OAI21_X1 _14966_ ( .A(\u_lsu.pmem[7140] ), .B1(_10880_ ), .B2(_11032_ ), .ZN(_11044_ ) );
AOI21_X1 _14967_ ( .A(fanout_net_20 ), .B1(_11043_ ), .B2(_11044_ ), .ZN(_00542_ ) );
NAND4_X1 _14968_ ( .A1(_10084_ ), .A2(_11042_ ), .A3(_11008_ ), .A4(_10997_ ), .ZN(_11045_ ) );
OAI21_X1 _14969_ ( .A(\u_lsu.pmem[7139] ), .B1(_10880_ ), .B2(_11032_ ), .ZN(_11046_ ) );
AOI21_X1 _14970_ ( .A(fanout_net_20 ), .B1(_11045_ ), .B2(_11046_ ), .ZN(_00543_ ) );
NAND4_X1 _14971_ ( .A1(_10088_ ), .A2(_11042_ ), .A3(_11008_ ), .A4(_10997_ ), .ZN(_11047_ ) );
BUF_X4 _14972_ ( .A(_10844_ ), .Z(_11048_ ) );
OAI21_X1 _14973_ ( .A(\u_lsu.pmem[7138] ), .B1(_11048_ ), .B2(_11032_ ), .ZN(_11049_ ) );
AOI21_X1 _14974_ ( .A(fanout_net_20 ), .B1(_11047_ ), .B2(_11049_ ), .ZN(_00544_ ) );
NAND4_X1 _14975_ ( .A1(_10094_ ), .A2(_11042_ ), .A3(_11008_ ), .A4(_10997_ ), .ZN(_11050_ ) );
OAI21_X1 _14976_ ( .A(\u_lsu.pmem[7137] ), .B1(_11048_ ), .B2(_11032_ ), .ZN(_11051_ ) );
AOI21_X1 _14977_ ( .A(fanout_net_20 ), .B1(_11050_ ), .B2(_11051_ ), .ZN(_00545_ ) );
NAND4_X1 _14978_ ( .A1(_10098_ ), .A2(_11042_ ), .A3(_11008_ ), .A4(_10997_ ), .ZN(_11052_ ) );
OAI21_X1 _14979_ ( .A(\u_lsu.pmem[7136] ), .B1(_11048_ ), .B2(_11032_ ), .ZN(_11053_ ) );
AOI21_X1 _14980_ ( .A(fanout_net_20 ), .B1(_11052_ ), .B2(_11053_ ), .ZN(_00546_ ) );
BUF_X4 _14981_ ( .A(_09572_ ), .Z(_11054_ ) );
INV_X1 _14982_ ( .A(_10102_ ), .ZN(_11055_ ) );
BUF_X4 _14983_ ( .A(_09664_ ), .Z(_11056_ ) );
NOR3_X1 _14984_ ( .A1(_10055_ ), .A2(_11055_ ), .A3(_11056_ ), .ZN(_11057_ ) );
NAND2_X1 _14985_ ( .A1(_11028_ ), .A2(_11057_ ), .ZN(_11058_ ) );
BUF_X4 _14986_ ( .A(_11058_ ), .Z(_11059_ ) );
OAI21_X1 _14987_ ( .A(\u_lsu.pmem[7111] ), .B1(_11054_ ), .B2(_11059_ ), .ZN(_11060_ ) );
BUF_X4 _14988_ ( .A(_10548_ ), .Z(_11061_ ) );
NAND4_X1 _14989_ ( .A1(_10851_ ), .A2(_11061_ ), .A3(_10993_ ), .A4(_11057_ ), .ZN(_11062_ ) );
AOI21_X1 _14990_ ( .A(fanout_net_21 ), .B1(_11060_ ), .B2(_11062_ ), .ZN(_00547_ ) );
BUF_X8 _14991_ ( .A(_09877_ ), .Z(_11063_ ) );
BUF_X4 _14992_ ( .A(_11063_ ), .Z(_11064_ ) );
NAND4_X1 _14993_ ( .A1(_10117_ ), .A2(_11042_ ), .A3(_11064_ ), .A4(_10997_ ), .ZN(_11065_ ) );
OAI21_X1 _14994_ ( .A(\u_lsu.pmem[7110] ), .B1(_11048_ ), .B2(_11059_ ), .ZN(_11066_ ) );
AOI21_X1 _14995_ ( .A(fanout_net_21 ), .B1(_11065_ ), .B2(_11066_ ), .ZN(_00548_ ) );
BUF_X4 _14996_ ( .A(_10592_ ), .Z(_11067_ ) );
NAND4_X1 _14997_ ( .A1(_10121_ ), .A2(_11042_ ), .A3(_11064_ ), .A4(_11067_ ), .ZN(_11068_ ) );
OAI21_X1 _14998_ ( .A(\u_lsu.pmem[7109] ), .B1(_11048_ ), .B2(_11059_ ), .ZN(_11069_ ) );
AOI21_X1 _14999_ ( .A(fanout_net_21 ), .B1(_11068_ ), .B2(_11069_ ), .ZN(_00549_ ) );
NAND4_X1 _15000_ ( .A1(_10125_ ), .A2(_11042_ ), .A3(_11064_ ), .A4(_11067_ ), .ZN(_11070_ ) );
OAI21_X1 _15001_ ( .A(\u_lsu.pmem[7108] ), .B1(_11048_ ), .B2(_11059_ ), .ZN(_11071_ ) );
AOI21_X1 _15002_ ( .A(fanout_net_21 ), .B1(_11070_ ), .B2(_11071_ ), .ZN(_00550_ ) );
NAND4_X1 _15003_ ( .A1(_10131_ ), .A2(_11042_ ), .A3(_11064_ ), .A4(_11067_ ), .ZN(_11072_ ) );
OAI21_X1 _15004_ ( .A(\u_lsu.pmem[7107] ), .B1(_11048_ ), .B2(_11059_ ), .ZN(_11073_ ) );
AOI21_X1 _15005_ ( .A(fanout_net_21 ), .B1(_11072_ ), .B2(_11073_ ), .ZN(_00551_ ) );
BUF_X4 _15006_ ( .A(_09675_ ), .Z(_11074_ ) );
NAND4_X1 _15007_ ( .A1(_10309_ ), .A2(_11039_ ), .A3(_11064_ ), .A4(_11074_ ), .ZN(_11075_ ) );
NAND2_X1 _15008_ ( .A1(_10944_ ), .A2(\u_lsu.pmem[3843] ), .ZN(_11076_ ) );
AOI21_X1 _15009_ ( .A(fanout_net_21 ), .B1(_11075_ ), .B2(_11076_ ), .ZN(_00552_ ) );
NAND4_X1 _15010_ ( .A1(_10135_ ), .A2(_11042_ ), .A3(_11064_ ), .A4(_11067_ ), .ZN(_11077_ ) );
OAI21_X1 _15011_ ( .A(\u_lsu.pmem[7106] ), .B1(_11048_ ), .B2(_11059_ ), .ZN(_11078_ ) );
AOI21_X1 _15012_ ( .A(fanout_net_21 ), .B1(_11077_ ), .B2(_11078_ ), .ZN(_00553_ ) );
BUF_X4 _15013_ ( .A(_09671_ ), .Z(_11079_ ) );
NAND4_X1 _15014_ ( .A1(_10138_ ), .A2(_11079_ ), .A3(_11064_ ), .A4(_11067_ ), .ZN(_11080_ ) );
OAI21_X1 _15015_ ( .A(\u_lsu.pmem[7105] ), .B1(_11048_ ), .B2(_11059_ ), .ZN(_11081_ ) );
AOI21_X1 _15016_ ( .A(fanout_net_21 ), .B1(_11080_ ), .B2(_11081_ ), .ZN(_00554_ ) );
NAND4_X1 _15017_ ( .A1(_10144_ ), .A2(_11079_ ), .A3(_11064_ ), .A4(_11067_ ), .ZN(_11082_ ) );
OAI21_X1 _15018_ ( .A(\u_lsu.pmem[7104] ), .B1(_11048_ ), .B2(_11059_ ), .ZN(_11083_ ) );
AOI21_X1 _15019_ ( .A(fanout_net_21 ), .B1(_11082_ ), .B2(_11083_ ), .ZN(_00555_ ) );
NAND4_X1 _15020_ ( .A1(_10148_ ), .A2(_11079_ ), .A3(_11064_ ), .A4(_11067_ ), .ZN(_11084_ ) );
BUF_X4 _15021_ ( .A(_10844_ ), .Z(_11085_ ) );
AND3_X2 _15022_ ( .A1(_09805_ ), .A2(_09784_ ), .A3(_09486_ ), .ZN(_11086_ ) );
NAND2_X1 _15023_ ( .A1(_11028_ ), .A2(_11086_ ), .ZN(_11087_ ) );
BUF_X4 _15024_ ( .A(_11087_ ), .Z(_11088_ ) );
OAI21_X1 _15025_ ( .A(\u_lsu.pmem[7079] ), .B1(_11085_ ), .B2(_11088_ ), .ZN(_11089_ ) );
AOI21_X1 _15026_ ( .A(fanout_net_21 ), .B1(_11084_ ), .B2(_11089_ ), .ZN(_00556_ ) );
NAND4_X1 _15027_ ( .A1(_10156_ ), .A2(_11079_ ), .A3(_11064_ ), .A4(_11067_ ), .ZN(_11090_ ) );
OAI21_X1 _15028_ ( .A(\u_lsu.pmem[7078] ), .B1(_11085_ ), .B2(_11088_ ), .ZN(_11091_ ) );
AOI21_X1 _15029_ ( .A(fanout_net_21 ), .B1(_11090_ ), .B2(_11091_ ), .ZN(_00557_ ) );
BUF_X4 _15030_ ( .A(_11063_ ), .Z(_11092_ ) );
NAND4_X1 _15031_ ( .A1(_10160_ ), .A2(_11079_ ), .A3(_11092_ ), .A4(_11067_ ), .ZN(_11093_ ) );
OAI21_X1 _15032_ ( .A(\u_lsu.pmem[7077] ), .B1(_11085_ ), .B2(_11088_ ), .ZN(_11094_ ) );
AOI21_X1 _15033_ ( .A(fanout_net_21 ), .B1(_11093_ ), .B2(_11094_ ), .ZN(_00558_ ) );
NAND4_X1 _15034_ ( .A1(_10166_ ), .A2(_11079_ ), .A3(_11092_ ), .A4(_11067_ ), .ZN(_11095_ ) );
OAI21_X1 _15035_ ( .A(\u_lsu.pmem[7076] ), .B1(_11085_ ), .B2(_11088_ ), .ZN(_11096_ ) );
AOI21_X1 _15036_ ( .A(fanout_net_21 ), .B1(_11095_ ), .B2(_11096_ ), .ZN(_00559_ ) );
BUF_X4 _15037_ ( .A(_10592_ ), .Z(_11097_ ) );
NAND4_X1 _15038_ ( .A1(_10169_ ), .A2(_11079_ ), .A3(_11092_ ), .A4(_11097_ ), .ZN(_11098_ ) );
OAI21_X1 _15039_ ( .A(\u_lsu.pmem[7075] ), .B1(_11085_ ), .B2(_11088_ ), .ZN(_11099_ ) );
AOI21_X1 _15040_ ( .A(fanout_net_21 ), .B1(_11098_ ), .B2(_11099_ ), .ZN(_00560_ ) );
NAND4_X1 _15041_ ( .A1(_10172_ ), .A2(_11079_ ), .A3(_11092_ ), .A4(_11097_ ), .ZN(_11100_ ) );
OAI21_X1 _15042_ ( .A(\u_lsu.pmem[7074] ), .B1(_11085_ ), .B2(_11088_ ), .ZN(_11101_ ) );
AOI21_X1 _15043_ ( .A(fanout_net_21 ), .B1(_11100_ ), .B2(_11101_ ), .ZN(_00561_ ) );
NAND4_X1 _15044_ ( .A1(_10176_ ), .A2(_11079_ ), .A3(_11092_ ), .A4(_11097_ ), .ZN(_11102_ ) );
OAI21_X1 _15045_ ( .A(\u_lsu.pmem[7073] ), .B1(_11085_ ), .B2(_11088_ ), .ZN(_11103_ ) );
AOI21_X1 _15046_ ( .A(fanout_net_21 ), .B1(_11102_ ), .B2(_11103_ ), .ZN(_00562_ ) );
NAND4_X1 _15047_ ( .A1(_10018_ ), .A2(_10887_ ), .A3(_11092_ ), .A4(_10313_ ), .ZN(_11104_ ) );
NAND2_X1 _15048_ ( .A1(_10944_ ), .A2(\u_lsu.pmem[3842] ), .ZN(_11105_ ) );
AOI21_X1 _15049_ ( .A(fanout_net_21 ), .B1(_11104_ ), .B2(_11105_ ), .ZN(_00563_ ) );
OAI21_X1 _15050_ ( .A(\u_lsu.pmem[7072] ), .B1(_11054_ ), .B2(_11088_ ), .ZN(_11106_ ) );
NAND4_X1 _15051_ ( .A1(_10525_ ), .A2(_11061_ ), .A3(_10993_ ), .A4(_11086_ ), .ZN(_11107_ ) );
AOI21_X1 _15052_ ( .A(fanout_net_21 ), .B1(_11106_ ), .B2(_11107_ ), .ZN(_00564_ ) );
AND3_X1 _15053_ ( .A1(_09504_ ), .A2(_09805_ ), .A3(_09462_ ), .ZN(_11108_ ) );
NAND2_X1 _15054_ ( .A1(_11108_ ), .A2(_11028_ ), .ZN(_11109_ ) );
BUF_X4 _15055_ ( .A(_11109_ ), .Z(_11110_ ) );
OAI21_X1 _15056_ ( .A(\u_lsu.pmem[7047] ), .B1(_11110_ ), .B2(_10936_ ), .ZN(_11111_ ) );
BUF_X4 _15057_ ( .A(_11108_ ), .Z(_11112_ ) );
BUF_X4 _15058_ ( .A(_11112_ ), .Z(_11113_ ) );
NAND4_X1 _15059_ ( .A1(_11113_ ), .A2(_10752_ ), .A3(_10993_ ), .A4(_10966_ ), .ZN(_11114_ ) );
AOI21_X1 _15060_ ( .A(fanout_net_21 ), .B1(_11111_ ), .B2(_11114_ ), .ZN(_00565_ ) );
OAI21_X1 _15061_ ( .A(\u_lsu.pmem[7046] ), .B1(_11110_ ), .B2(_10936_ ), .ZN(_11115_ ) );
NAND4_X1 _15062_ ( .A1(_11113_ ), .A2(_10185_ ), .A3(_10993_ ), .A4(_10966_ ), .ZN(_11116_ ) );
AOI21_X1 _15063_ ( .A(fanout_net_21 ), .B1(_11115_ ), .B2(_11116_ ), .ZN(_00566_ ) );
OAI21_X1 _15064_ ( .A(\u_lsu.pmem[7045] ), .B1(_11110_ ), .B2(_10936_ ), .ZN(_11117_ ) );
NAND4_X1 _15065_ ( .A1(_11113_ ), .A2(_10188_ ), .A3(_10993_ ), .A4(_10966_ ), .ZN(_11118_ ) );
AOI21_X1 _15066_ ( .A(fanout_net_21 ), .B1(_11117_ ), .B2(_11118_ ), .ZN(_00567_ ) );
OAI21_X1 _15067_ ( .A(\u_lsu.pmem[7044] ), .B1(_11110_ ), .B2(_10936_ ), .ZN(_11119_ ) );
NAND4_X1 _15068_ ( .A1(_11113_ ), .A2(_10192_ ), .A3(_10993_ ), .A4(_10966_ ), .ZN(_11120_ ) );
AOI21_X1 _15069_ ( .A(fanout_net_21 ), .B1(_11119_ ), .B2(_11120_ ), .ZN(_00568_ ) );
OAI21_X1 _15070_ ( .A(\u_lsu.pmem[7043] ), .B1(_11110_ ), .B2(_10936_ ), .ZN(_11121_ ) );
NAND4_X1 _15071_ ( .A1(_11113_ ), .A2(_10915_ ), .A3(_10993_ ), .A4(_10966_ ), .ZN(_11122_ ) );
AOI21_X1 _15072_ ( .A(fanout_net_21 ), .B1(_11121_ ), .B2(_11122_ ), .ZN(_00569_ ) );
BUF_X4 _15073_ ( .A(_10901_ ), .Z(_11123_ ) );
OAI21_X1 _15074_ ( .A(\u_lsu.pmem[7042] ), .B1(_11110_ ), .B2(_11123_ ), .ZN(_11124_ ) );
BUF_X4 _15075_ ( .A(_09878_ ), .Z(_11125_ ) );
NAND4_X1 _15076_ ( .A1(_09874_ ), .A2(_09540_ ), .A3(_11125_ ), .A4(_10966_ ), .ZN(_11126_ ) );
AOI21_X1 _15077_ ( .A(fanout_net_21 ), .B1(_11124_ ), .B2(_11126_ ), .ZN(_00570_ ) );
OAI21_X1 _15078_ ( .A(\u_lsu.pmem[7041] ), .B1(_11110_ ), .B2(_11123_ ), .ZN(_11127_ ) );
BUF_X4 _15079_ ( .A(_10904_ ), .Z(_11128_ ) );
NAND4_X1 _15080_ ( .A1(_11113_ ), .A2(_09923_ ), .A3(_11125_ ), .A4(_11128_ ), .ZN(_11129_ ) );
AOI21_X1 _15081_ ( .A(fanout_net_21 ), .B1(_11127_ ), .B2(_11129_ ), .ZN(_00571_ ) );
OAI21_X1 _15082_ ( .A(\u_lsu.pmem[7040] ), .B1(_11110_ ), .B2(_11123_ ), .ZN(_11130_ ) );
BUF_X4 _15083_ ( .A(_09547_ ), .Z(_11131_ ) );
NAND4_X1 _15084_ ( .A1(_11113_ ), .A2(_11131_ ), .A3(_11125_ ), .A4(_11128_ ), .ZN(_11132_ ) );
AOI21_X1 _15085_ ( .A(fanout_net_21 ), .B1(_11130_ ), .B2(_11132_ ), .ZN(_00572_ ) );
AND2_X1 _15086_ ( .A1(_10008_ ), .A2(_08995_ ), .ZN(_11133_ ) );
AND2_X2 _15087_ ( .A1(_10325_ ), .A2(_11133_ ), .ZN(_11134_ ) );
INV_X1 _15088_ ( .A(_11134_ ), .ZN(_11135_ ) );
BUF_X4 _15089_ ( .A(_11135_ ), .Z(_11136_ ) );
OAI21_X1 _15090_ ( .A(\u_lsu.pmem[7015] ), .B1(_11054_ ), .B2(_11136_ ), .ZN(_11137_ ) );
BUF_X4 _15091_ ( .A(_09741_ ), .Z(_11138_ ) );
BUF_X4 _15092_ ( .A(_09635_ ), .Z(_11139_ ) );
BUF_X4 _15093_ ( .A(_11134_ ), .Z(_11140_ ) );
NAND3_X1 _15094_ ( .A1(_11138_ ), .A2(_11139_ ), .A3(_11140_ ), .ZN(_11141_ ) );
AOI21_X1 _15095_ ( .A(fanout_net_21 ), .B1(_11137_ ), .B2(_11141_ ), .ZN(_00573_ ) );
NAND4_X1 _15096_ ( .A1(_10316_ ), .A2(_11039_ ), .A3(_11092_ ), .A4(_11074_ ), .ZN(_11142_ ) );
NAND2_X1 _15097_ ( .A1(_10944_ ), .A2(\u_lsu.pmem[3841] ), .ZN(_11143_ ) );
AOI21_X1 _15098_ ( .A(fanout_net_21 ), .B1(_11142_ ), .B2(_11143_ ), .ZN(_00574_ ) );
OAI21_X1 _15099_ ( .A(\u_lsu.pmem[7014] ), .B1(_11054_ ), .B2(_11136_ ), .ZN(_11144_ ) );
BUF_X4 _15100_ ( .A(_09578_ ), .Z(_11145_ ) );
NAND3_X1 _15101_ ( .A1(_11145_ ), .A2(_11139_ ), .A3(_11140_ ), .ZN(_11146_ ) );
AOI21_X1 _15102_ ( .A(fanout_net_21 ), .B1(_11144_ ), .B2(_11146_ ), .ZN(_00575_ ) );
OAI21_X1 _15103_ ( .A(\u_lsu.pmem[7013] ), .B1(_11054_ ), .B2(_11135_ ), .ZN(_11147_ ) );
BUF_X4 _15104_ ( .A(_09585_ ), .Z(_11148_ ) );
NAND3_X1 _15105_ ( .A1(_11148_ ), .A2(_11139_ ), .A3(_11140_ ), .ZN(_11149_ ) );
AOI21_X1 _15106_ ( .A(fanout_net_21 ), .B1(_11147_ ), .B2(_11149_ ), .ZN(_00576_ ) );
OAI21_X1 _15107_ ( .A(\u_lsu.pmem[7012] ), .B1(_11054_ ), .B2(_11135_ ), .ZN(_11150_ ) );
BUF_X4 _15108_ ( .A(_09147_ ), .Z(_11151_ ) );
BUF_X4 _15109_ ( .A(_11151_ ), .Z(_11152_ ) );
NAND3_X1 _15110_ ( .A1(_11152_ ), .A2(_11139_ ), .A3(_11140_ ), .ZN(_11153_ ) );
AOI21_X1 _15111_ ( .A(fanout_net_22 ), .B1(_11150_ ), .B2(_11153_ ), .ZN(_00577_ ) );
OAI21_X1 _15112_ ( .A(\u_lsu.pmem[7011] ), .B1(_11054_ ), .B2(_11135_ ), .ZN(_11154_ ) );
BUF_X4 _15113_ ( .A(_09448_ ), .Z(_11155_ ) );
NAND3_X1 _15114_ ( .A1(_11155_ ), .A2(_11139_ ), .A3(_11140_ ), .ZN(_11156_ ) );
AOI21_X1 _15115_ ( .A(fanout_net_22 ), .B1(_11154_ ), .B2(_11156_ ), .ZN(_00578_ ) );
OAI21_X1 _15116_ ( .A(\u_lsu.pmem[7010] ), .B1(_11054_ ), .B2(_11135_ ), .ZN(_11157_ ) );
BUF_X4 _15117_ ( .A(_09611_ ), .Z(_11158_ ) );
BUF_X4 _15118_ ( .A(_09141_ ), .Z(_11159_ ) );
BUF_X4 _15119_ ( .A(_11159_ ), .Z(_11160_ ) );
NAND3_X1 _15120_ ( .A1(_11158_ ), .A2(_11160_ ), .A3(_11140_ ), .ZN(_11161_ ) );
AOI21_X1 _15121_ ( .A(fanout_net_22 ), .B1(_11157_ ), .B2(_11161_ ), .ZN(_00579_ ) );
OAI21_X1 _15122_ ( .A(\u_lsu.pmem[7009] ), .B1(_11054_ ), .B2(_11135_ ), .ZN(_11162_ ) );
BUF_X4 _15123_ ( .A(_09616_ ), .Z(_11163_ ) );
NAND3_X1 _15124_ ( .A1(_11163_ ), .A2(_11160_ ), .A3(_11140_ ), .ZN(_11164_ ) );
AOI21_X1 _15125_ ( .A(fanout_net_22 ), .B1(_11162_ ), .B2(_11164_ ), .ZN(_00580_ ) );
OAI21_X1 _15126_ ( .A(\u_lsu.pmem[7008] ), .B1(_11054_ ), .B2(_11135_ ), .ZN(_11165_ ) );
NAND3_X1 _15127_ ( .A1(_10741_ ), .A2(_11160_ ), .A3(_11140_ ), .ZN(_11166_ ) );
AOI21_X1 _15128_ ( .A(fanout_net_22 ), .B1(_11165_ ), .B2(_11166_ ), .ZN(_00581_ ) );
BUF_X4 _15129_ ( .A(_09572_ ), .Z(_11167_ ) );
AND2_X1 _15130_ ( .A1(_10226_ ), .A2(_08995_ ), .ZN(_11168_ ) );
AND2_X2 _15131_ ( .A1(_10325_ ), .A2(_11168_ ), .ZN(_11169_ ) );
INV_X1 _15132_ ( .A(_11169_ ), .ZN(_11170_ ) );
BUF_X4 _15133_ ( .A(_11170_ ), .Z(_11171_ ) );
OAI21_X1 _15134_ ( .A(\u_lsu.pmem[6983] ), .B1(_11167_ ), .B2(_11171_ ), .ZN(_11172_ ) );
BUF_X4 _15135_ ( .A(_11169_ ), .Z(_11173_ ) );
NAND3_X1 _15136_ ( .A1(_11138_ ), .A2(_11160_ ), .A3(_11173_ ), .ZN(_11174_ ) );
AOI21_X1 _15137_ ( .A(fanout_net_22 ), .B1(_11172_ ), .B2(_11174_ ), .ZN(_00582_ ) );
OAI21_X1 _15138_ ( .A(\u_lsu.pmem[6982] ), .B1(_11167_ ), .B2(_11171_ ), .ZN(_11175_ ) );
NAND3_X1 _15139_ ( .A1(_10719_ ), .A2(_11160_ ), .A3(_11173_ ), .ZN(_11176_ ) );
AOI21_X1 _15140_ ( .A(fanout_net_22 ), .B1(_11175_ ), .B2(_11176_ ), .ZN(_00583_ ) );
OAI21_X1 _15141_ ( .A(\u_lsu.pmem[6981] ), .B1(_11167_ ), .B2(_11170_ ), .ZN(_11177_ ) );
NAND3_X1 _15142_ ( .A1(_10728_ ), .A2(_11160_ ), .A3(_11173_ ), .ZN(_11178_ ) );
AOI21_X1 _15143_ ( .A(fanout_net_22 ), .B1(_11177_ ), .B2(_11178_ ), .ZN(_00584_ ) );
NAND4_X1 _15144_ ( .A1(_09756_ ), .A2(_11079_ ), .A3(_09869_ ), .A4(_11097_ ), .ZN(_11179_ ) );
OAI21_X1 _15145_ ( .A(\u_lsu.pmem[4326] ), .B1(_11085_ ), .B2(_09752_ ), .ZN(_11180_ ) );
AOI21_X1 _15146_ ( .A(fanout_net_22 ), .B1(_11179_ ), .B2(_11180_ ), .ZN(_00585_ ) );
NAND4_X1 _15147_ ( .A1(_10320_ ), .A2(_11039_ ), .A3(_11092_ ), .A4(_11074_ ), .ZN(_11181_ ) );
NAND2_X1 _15148_ ( .A1(_10944_ ), .A2(\u_lsu.pmem[3840] ), .ZN(_11182_ ) );
AOI21_X1 _15149_ ( .A(fanout_net_22 ), .B1(_11181_ ), .B2(_11182_ ), .ZN(_00586_ ) );
OAI21_X1 _15150_ ( .A(\u_lsu.pmem[6980] ), .B1(_11167_ ), .B2(_11170_ ), .ZN(_11183_ ) );
NAND3_X1 _15151_ ( .A1(_11152_ ), .A2(_11160_ ), .A3(_11173_ ), .ZN(_11184_ ) );
AOI21_X1 _15152_ ( .A(fanout_net_22 ), .B1(_11183_ ), .B2(_11184_ ), .ZN(_00587_ ) );
OAI21_X1 _15153_ ( .A(\u_lsu.pmem[6979] ), .B1(_11167_ ), .B2(_11170_ ), .ZN(_11185_ ) );
NAND3_X1 _15154_ ( .A1(_11155_ ), .A2(_11160_ ), .A3(_11173_ ), .ZN(_11186_ ) );
AOI21_X1 _15155_ ( .A(fanout_net_22 ), .B1(_11185_ ), .B2(_11186_ ), .ZN(_00588_ ) );
OAI21_X1 _15156_ ( .A(\u_lsu.pmem[6978] ), .B1(_11167_ ), .B2(_11170_ ), .ZN(_11187_ ) );
NAND3_X1 _15157_ ( .A1(_11158_ ), .A2(_11160_ ), .A3(_11173_ ), .ZN(_11188_ ) );
AOI21_X1 _15158_ ( .A(fanout_net_22 ), .B1(_11187_ ), .B2(_11188_ ), .ZN(_00589_ ) );
OAI21_X1 _15159_ ( .A(\u_lsu.pmem[6977] ), .B1(_11167_ ), .B2(_11170_ ), .ZN(_11189_ ) );
NAND3_X1 _15160_ ( .A1(_11163_ ), .A2(_11160_ ), .A3(_11173_ ), .ZN(_11190_ ) );
AOI21_X1 _15161_ ( .A(fanout_net_22 ), .B1(_11189_ ), .B2(_11190_ ), .ZN(_00590_ ) );
OAI21_X1 _15162_ ( .A(\u_lsu.pmem[6976] ), .B1(_11167_ ), .B2(_11170_ ), .ZN(_11191_ ) );
BUF_X4 _15163_ ( .A(_09635_ ), .Z(_11192_ ) );
NAND3_X1 _15164_ ( .A1(_10741_ ), .A2(_11192_ ), .A3(_11173_ ), .ZN(_11193_ ) );
AOI21_X1 _15165_ ( .A(fanout_net_22 ), .B1(_11191_ ), .B2(_11193_ ), .ZN(_00591_ ) );
BUF_X4 _15166_ ( .A(_09671_ ), .Z(_11194_ ) );
NAND4_X1 _15167_ ( .A1(_10250_ ), .A2(_11194_ ), .A3(_11092_ ), .A4(_11097_ ), .ZN(_11195_ ) );
BUF_X4 _15168_ ( .A(_09664_ ), .Z(_11196_ ) );
NOR3_X1 _15169_ ( .A1(_10009_ ), .A2(_09128_ ), .A3(_11196_ ), .ZN(_11197_ ) );
AND2_X2 _15170_ ( .A1(_09135_ ), .A2(_11197_ ), .ZN(_11198_ ) );
INV_X1 _15171_ ( .A(_11198_ ), .ZN(_11199_ ) );
OAI21_X1 _15172_ ( .A(\u_lsu.pmem[6951] ), .B1(_11085_ ), .B2(_11199_ ), .ZN(_11200_ ) );
AOI21_X1 _15173_ ( .A(fanout_net_22 ), .B1(_11195_ ), .B2(_11200_ ), .ZN(_00592_ ) );
NAND4_X1 _15174_ ( .A1(_10263_ ), .A2(_11194_ ), .A3(_11092_ ), .A4(_11097_ ), .ZN(_11201_ ) );
OAI21_X1 _15175_ ( .A(\u_lsu.pmem[6950] ), .B1(_11085_ ), .B2(_11199_ ), .ZN(_11202_ ) );
AOI21_X1 _15176_ ( .A(fanout_net_22 ), .B1(_11201_ ), .B2(_11202_ ), .ZN(_00593_ ) );
BUF_X4 _15177_ ( .A(_11063_ ), .Z(_11203_ ) );
NAND4_X1 _15178_ ( .A1(_10267_ ), .A2(_11194_ ), .A3(_11203_ ), .A4(_11097_ ), .ZN(_11204_ ) );
BUF_X4 _15179_ ( .A(_10844_ ), .Z(_11205_ ) );
OAI21_X1 _15180_ ( .A(\u_lsu.pmem[6949] ), .B1(_11205_ ), .B2(_11199_ ), .ZN(_11206_ ) );
AOI21_X1 _15181_ ( .A(fanout_net_22 ), .B1(_11204_ ), .B2(_11206_ ), .ZN(_00594_ ) );
AND2_X1 _15182_ ( .A1(_09141_ ), .A2(_11198_ ), .ZN(_11207_ ) );
OAI21_X1 _15183_ ( .A(_10715_ ), .B1(_11207_ ), .B2(\u_lsu.pmem[6948] ), .ZN(_11208_ ) );
AOI21_X1 _15184_ ( .A(_11208_ ), .B1(_09691_ ), .B2(_11207_ ), .ZN(_00595_ ) );
BUF_X4 _15185_ ( .A(_11199_ ), .Z(_11209_ ) );
OAI21_X1 _15186_ ( .A(\u_lsu.pmem[6947] ), .B1(_11167_ ), .B2(_11209_ ), .ZN(_11210_ ) );
NAND3_X1 _15187_ ( .A1(_11155_ ), .A2(_11192_ ), .A3(_11198_ ), .ZN(_11211_ ) );
AOI21_X1 _15188_ ( .A(fanout_net_22 ), .B1(_11210_ ), .B2(_11211_ ), .ZN(_00596_ ) );
BUF_X4 _15189_ ( .A(_10065_ ), .Z(_11212_ ) );
NAND4_X1 _15190_ ( .A1(_10018_ ), .A2(_11212_ ), .A3(_09914_ ), .A4(_10324_ ), .ZN(_11213_ ) );
BUF_X4 _15191_ ( .A(_09472_ ), .Z(_11214_ ) );
OAI21_X1 _15192_ ( .A(\u_lsu.pmem[3815] ), .B1(_11214_ ), .B2(_10328_ ), .ZN(_11215_ ) );
AOI21_X1 _15193_ ( .A(fanout_net_22 ), .B1(_11213_ ), .B2(_11215_ ), .ZN(_00597_ ) );
OAI21_X1 _15194_ ( .A(\u_lsu.pmem[6946] ), .B1(_11167_ ), .B2(_11209_ ), .ZN(_11216_ ) );
NAND3_X1 _15195_ ( .A1(_11158_ ), .A2(_11192_ ), .A3(_11198_ ), .ZN(_11217_ ) );
AOI21_X1 _15196_ ( .A(fanout_net_22 ), .B1(_11216_ ), .B2(_11217_ ), .ZN(_00598_ ) );
BUF_X4 _15197_ ( .A(_09572_ ), .Z(_11218_ ) );
OAI21_X1 _15198_ ( .A(\u_lsu.pmem[6945] ), .B1(_11218_ ), .B2(_11209_ ), .ZN(_11219_ ) );
NAND3_X1 _15199_ ( .A1(_11163_ ), .A2(_11192_ ), .A3(_11198_ ), .ZN(_11220_ ) );
AOI21_X1 _15200_ ( .A(fanout_net_22 ), .B1(_11219_ ), .B2(_11220_ ), .ZN(_00599_ ) );
NAND4_X1 _15201_ ( .A1(_10279_ ), .A2(_11194_ ), .A3(_11203_ ), .A4(_11097_ ), .ZN(_11221_ ) );
OAI21_X1 _15202_ ( .A(\u_lsu.pmem[6944] ), .B1(_11205_ ), .B2(_11199_ ), .ZN(_11222_ ) );
AOI21_X1 _15203_ ( .A(fanout_net_22 ), .B1(_11221_ ), .B2(_11222_ ), .ZN(_00600_ ) );
NAND4_X1 _15204_ ( .A1(_10285_ ), .A2(_11194_ ), .A3(_11203_ ), .A4(_11097_ ), .ZN(_11223_ ) );
NAND3_X1 _15205_ ( .A1(_10424_ ), .A2(_09842_ ), .A3(_10289_ ), .ZN(_11224_ ) );
BUF_X4 _15206_ ( .A(_11224_ ), .Z(_11225_ ) );
OAI21_X1 _15207_ ( .A(\u_lsu.pmem[6919] ), .B1(_11205_ ), .B2(_11225_ ), .ZN(_11226_ ) );
AOI21_X1 _15208_ ( .A(fanout_net_22 ), .B1(_11223_ ), .B2(_11226_ ), .ZN(_00601_ ) );
NAND4_X1 _15209_ ( .A1(_10295_ ), .A2(_11194_ ), .A3(_11203_ ), .A4(_11097_ ), .ZN(_11227_ ) );
OAI21_X1 _15210_ ( .A(\u_lsu.pmem[6918] ), .B1(_11205_ ), .B2(_11225_ ), .ZN(_11228_ ) );
AOI21_X1 _15211_ ( .A(fanout_net_22 ), .B1(_11227_ ), .B2(_11228_ ), .ZN(_00602_ ) );
BUF_X4 _15212_ ( .A(_10592_ ), .Z(_11229_ ) );
NAND4_X1 _15213_ ( .A1(_10299_ ), .A2(_11194_ ), .A3(_11203_ ), .A4(_11229_ ), .ZN(_11230_ ) );
OAI21_X1 _15214_ ( .A(\u_lsu.pmem[6917] ), .B1(_11205_ ), .B2(_11225_ ), .ZN(_11231_ ) );
AOI21_X1 _15215_ ( .A(fanout_net_22 ), .B1(_11230_ ), .B2(_11231_ ), .ZN(_00603_ ) );
NAND4_X1 _15216_ ( .A1(_10306_ ), .A2(_11194_ ), .A3(_11203_ ), .A4(_11229_ ), .ZN(_11232_ ) );
OAI21_X1 _15217_ ( .A(\u_lsu.pmem[6916] ), .B1(_11205_ ), .B2(_11225_ ), .ZN(_11233_ ) );
AOI21_X1 _15218_ ( .A(fanout_net_22 ), .B1(_11232_ ), .B2(_11233_ ), .ZN(_00604_ ) );
NAND4_X1 _15219_ ( .A1(_10309_ ), .A2(_11194_ ), .A3(_11203_ ), .A4(_11229_ ), .ZN(_11234_ ) );
OAI21_X1 _15220_ ( .A(\u_lsu.pmem[6915] ), .B1(_11205_ ), .B2(_11225_ ), .ZN(_11235_ ) );
AOI21_X1 _15221_ ( .A(fanout_net_22 ), .B1(_11234_ ), .B2(_11235_ ), .ZN(_00605_ ) );
OAI21_X1 _15222_ ( .A(\u_lsu.pmem[6914] ), .B1(_11218_ ), .B2(_11225_ ), .ZN(_11236_ ) );
NAND4_X1 _15223_ ( .A1(_09510_ ), .A2(_09540_ ), .A3(_11125_ ), .A4(_10313_ ), .ZN(_11237_ ) );
AOI21_X1 _15224_ ( .A(fanout_net_22 ), .B1(_11236_ ), .B2(_11237_ ), .ZN(_00606_ ) );
NAND4_X1 _15225_ ( .A1(_10316_ ), .A2(_11194_ ), .A3(_11203_ ), .A4(_11229_ ), .ZN(_11238_ ) );
OAI21_X1 _15226_ ( .A(\u_lsu.pmem[6913] ), .B1(_11205_ ), .B2(_11225_ ), .ZN(_11239_ ) );
AOI21_X1 _15227_ ( .A(fanout_net_22 ), .B1(_11238_ ), .B2(_11239_ ), .ZN(_00607_ ) );
NAND4_X1 _15228_ ( .A1(_10332_ ), .A2(_10887_ ), .A3(_11203_ ), .A4(_11074_ ), .ZN(_11240_ ) );
OAI21_X1 _15229_ ( .A(\u_lsu.pmem[3814] ), .B1(_11214_ ), .B2(_10328_ ), .ZN(_11241_ ) );
AOI21_X1 _15230_ ( .A(fanout_net_23 ), .B1(_11240_ ), .B2(_11241_ ), .ZN(_00608_ ) );
BUF_X4 _15231_ ( .A(_09671_ ), .Z(_11242_ ) );
NAND4_X1 _15232_ ( .A1(_10320_ ), .A2(_11242_ ), .A3(_11203_ ), .A4(_11229_ ), .ZN(_11243_ ) );
OAI21_X1 _15233_ ( .A(\u_lsu.pmem[6912] ), .B1(_11205_ ), .B2(_11225_ ), .ZN(_11244_ ) );
AOI21_X1 _15234_ ( .A(fanout_net_23 ), .B1(_11243_ ), .B2(_11244_ ), .ZN(_00609_ ) );
NOR2_X1 _15235_ ( .A1(_10323_ ), .A2(_10397_ ), .ZN(_11245_ ) );
NAND2_X1 _15236_ ( .A1(_11245_ ), .A2(_10424_ ), .ZN(_11246_ ) );
BUF_X4 _15237_ ( .A(_11246_ ), .Z(_11247_ ) );
OAI21_X1 _15238_ ( .A(\u_lsu.pmem[6887] ), .B1(_11218_ ), .B2(_11247_ ), .ZN(_11248_ ) );
NAND4_X1 _15239_ ( .A1(_10851_ ), .A2(_11061_ ), .A3(_11125_ ), .A4(_11245_ ), .ZN(_11249_ ) );
AOI21_X1 _15240_ ( .A(fanout_net_23 ), .B1(_11248_ ), .B2(_11249_ ), .ZN(_00610_ ) );
BUF_X4 _15241_ ( .A(_11063_ ), .Z(_11250_ ) );
NAND4_X1 _15242_ ( .A1(_10332_ ), .A2(_11242_ ), .A3(_11250_ ), .A4(_11229_ ), .ZN(_11251_ ) );
OAI21_X1 _15243_ ( .A(\u_lsu.pmem[6886] ), .B1(_11205_ ), .B2(_11247_ ), .ZN(_11252_ ) );
AOI21_X1 _15244_ ( .A(fanout_net_23 ), .B1(_11251_ ), .B2(_11252_ ), .ZN(_00611_ ) );
NAND4_X1 _15245_ ( .A1(_10336_ ), .A2(_11242_ ), .A3(_11250_ ), .A4(_11229_ ), .ZN(_11253_ ) );
BUF_X4 _15246_ ( .A(_10844_ ), .Z(_11254_ ) );
OAI21_X1 _15247_ ( .A(\u_lsu.pmem[6885] ), .B1(_11254_ ), .B2(_11247_ ), .ZN(_11255_ ) );
AOI21_X1 _15248_ ( .A(fanout_net_23 ), .B1(_11253_ ), .B2(_11255_ ), .ZN(_00612_ ) );
NAND4_X1 _15249_ ( .A1(_10339_ ), .A2(_11242_ ), .A3(_11250_ ), .A4(_11229_ ), .ZN(_11256_ ) );
OAI21_X1 _15250_ ( .A(\u_lsu.pmem[6884] ), .B1(_11254_ ), .B2(_11247_ ), .ZN(_11257_ ) );
AOI21_X1 _15251_ ( .A(fanout_net_23 ), .B1(_11256_ ), .B2(_11257_ ), .ZN(_00613_ ) );
NAND4_X1 _15252_ ( .A1(_10345_ ), .A2(_11242_ ), .A3(_11250_ ), .A4(_11229_ ), .ZN(_11258_ ) );
OAI21_X1 _15253_ ( .A(\u_lsu.pmem[6883] ), .B1(_11254_ ), .B2(_11247_ ), .ZN(_11259_ ) );
AOI21_X1 _15254_ ( .A(fanout_net_23 ), .B1(_11258_ ), .B2(_11259_ ), .ZN(_00614_ ) );
NAND4_X1 _15255_ ( .A1(_10350_ ), .A2(_11242_ ), .A3(_11250_ ), .A4(_11229_ ), .ZN(_11260_ ) );
OAI21_X1 _15256_ ( .A(\u_lsu.pmem[6882] ), .B1(_11254_ ), .B2(_11247_ ), .ZN(_11261_ ) );
AOI21_X1 _15257_ ( .A(fanout_net_23 ), .B1(_11260_ ), .B2(_11261_ ), .ZN(_00615_ ) );
BUF_X4 _15258_ ( .A(_10592_ ), .Z(_11262_ ) );
NAND4_X1 _15259_ ( .A1(_10354_ ), .A2(_11242_ ), .A3(_11250_ ), .A4(_11262_ ), .ZN(_11263_ ) );
OAI21_X1 _15260_ ( .A(\u_lsu.pmem[6881] ), .B1(_11254_ ), .B2(_11247_ ), .ZN(_11264_ ) );
AOI21_X1 _15261_ ( .A(fanout_net_23 ), .B1(_11263_ ), .B2(_11264_ ), .ZN(_00616_ ) );
NAND4_X1 _15262_ ( .A1(_10357_ ), .A2(_11242_ ), .A3(_11250_ ), .A4(_11262_ ), .ZN(_11265_ ) );
OAI21_X1 _15263_ ( .A(\u_lsu.pmem[6880] ), .B1(_11254_ ), .B2(_11247_ ), .ZN(_11266_ ) );
AOI21_X1 _15264_ ( .A(fanout_net_23 ), .B1(_11265_ ), .B2(_11266_ ), .ZN(_00617_ ) );
NOR2_X1 _15265_ ( .A1(_10361_ ), .A2(_10397_ ), .ZN(_11267_ ) );
NAND2_X1 _15266_ ( .A1(_11267_ ), .A2(_10424_ ), .ZN(_11268_ ) );
BUF_X4 _15267_ ( .A(_11268_ ), .Z(_11269_ ) );
OAI21_X1 _15268_ ( .A(\u_lsu.pmem[6855] ), .B1(_11218_ ), .B2(_11269_ ), .ZN(_11270_ ) );
NAND4_X1 _15269_ ( .A1(_10851_ ), .A2(_11061_ ), .A3(_11125_ ), .A4(_11267_ ), .ZN(_11271_ ) );
AOI21_X1 _15270_ ( .A(fanout_net_23 ), .B1(_11270_ ), .B2(_11271_ ), .ZN(_00618_ ) );
NAND4_X1 _15271_ ( .A1(_10336_ ), .A2(_10887_ ), .A3(_11250_ ), .A4(_11074_ ), .ZN(_11272_ ) );
OAI21_X1 _15272_ ( .A(\u_lsu.pmem[3813] ), .B1(_11214_ ), .B2(_10327_ ), .ZN(_11273_ ) );
AOI21_X1 _15273_ ( .A(fanout_net_23 ), .B1(_11272_ ), .B2(_11273_ ), .ZN(_00619_ ) );
NAND4_X1 _15274_ ( .A1(_10368_ ), .A2(_11242_ ), .A3(_11250_ ), .A4(_11262_ ), .ZN(_11274_ ) );
OAI21_X1 _15275_ ( .A(\u_lsu.pmem[6854] ), .B1(_11254_ ), .B2(_11269_ ), .ZN(_11275_ ) );
AOI21_X1 _15276_ ( .A(fanout_net_23 ), .B1(_11274_ ), .B2(_11275_ ), .ZN(_00620_ ) );
NAND4_X1 _15277_ ( .A1(_10371_ ), .A2(_11242_ ), .A3(_11250_ ), .A4(_11262_ ), .ZN(_11276_ ) );
OAI21_X1 _15278_ ( .A(\u_lsu.pmem[6853] ), .B1(_11254_ ), .B2(_11269_ ), .ZN(_11277_ ) );
AOI21_X1 _15279_ ( .A(fanout_net_23 ), .B1(_11276_ ), .B2(_11277_ ), .ZN(_00621_ ) );
BUF_X4 _15280_ ( .A(_09671_ ), .Z(_11278_ ) );
BUF_X4 _15281_ ( .A(_11063_ ), .Z(_11279_ ) );
NAND4_X1 _15282_ ( .A1(_10374_ ), .A2(_11278_ ), .A3(_11279_ ), .A4(_11262_ ), .ZN(_11280_ ) );
OAI21_X1 _15283_ ( .A(\u_lsu.pmem[6852] ), .B1(_11254_ ), .B2(_11269_ ), .ZN(_11281_ ) );
AOI21_X1 _15284_ ( .A(fanout_net_23 ), .B1(_11280_ ), .B2(_11281_ ), .ZN(_00622_ ) );
NAND4_X1 _15285_ ( .A1(_10377_ ), .A2(_11278_ ), .A3(_11279_ ), .A4(_11262_ ), .ZN(_11282_ ) );
OAI21_X1 _15286_ ( .A(\u_lsu.pmem[6851] ), .B1(_11254_ ), .B2(_11269_ ), .ZN(_11283_ ) );
AOI21_X1 _15287_ ( .A(fanout_net_23 ), .B1(_11282_ ), .B2(_11283_ ), .ZN(_00623_ ) );
NAND4_X1 _15288_ ( .A1(_10381_ ), .A2(_11278_ ), .A3(_11279_ ), .A4(_11262_ ), .ZN(_11284_ ) );
BUF_X4 _15289_ ( .A(_10844_ ), .Z(_11285_ ) );
OAI21_X1 _15290_ ( .A(\u_lsu.pmem[6850] ), .B1(_11285_ ), .B2(_11269_ ), .ZN(_11286_ ) );
AOI21_X1 _15291_ ( .A(fanout_net_23 ), .B1(_11284_ ), .B2(_11286_ ), .ZN(_00624_ ) );
NAND4_X1 _15292_ ( .A1(_10384_ ), .A2(_11278_ ), .A3(_11279_ ), .A4(_11262_ ), .ZN(_11287_ ) );
OAI21_X1 _15293_ ( .A(\u_lsu.pmem[6849] ), .B1(_11285_ ), .B2(_11269_ ), .ZN(_11288_ ) );
AOI21_X1 _15294_ ( .A(fanout_net_23 ), .B1(_11287_ ), .B2(_11288_ ), .ZN(_00625_ ) );
NAND4_X1 _15295_ ( .A1(_10391_ ), .A2(_11278_ ), .A3(_11279_ ), .A4(_11262_ ), .ZN(_11289_ ) );
OAI21_X1 _15296_ ( .A(\u_lsu.pmem[6848] ), .B1(_11285_ ), .B2(_11269_ ), .ZN(_11290_ ) );
AOI21_X1 _15297_ ( .A(fanout_net_23 ), .B1(_11289_ ), .B2(_11290_ ), .ZN(_00626_ ) );
NAND4_X1 _15298_ ( .A1(_10394_ ), .A2(_11278_ ), .A3(_11279_ ), .A4(_11262_ ), .ZN(_11291_ ) );
AND3_X2 _15299_ ( .A1(_09538_ ), .A2(_09462_ ), .A3(_09857_ ), .ZN(_11292_ ) );
NAND2_X1 _15300_ ( .A1(_11292_ ), .A2(_11028_ ), .ZN(_11293_ ) );
BUF_X4 _15301_ ( .A(_11293_ ), .Z(_11294_ ) );
OAI21_X1 _15302_ ( .A(\u_lsu.pmem[6823] ), .B1(_11285_ ), .B2(_11294_ ), .ZN(_11295_ ) );
AOI21_X1 _15303_ ( .A(fanout_net_23 ), .B1(_11291_ ), .B2(_11295_ ), .ZN(_00627_ ) );
BUF_X4 _15304_ ( .A(_10592_ ), .Z(_11296_ ) );
NAND4_X1 _15305_ ( .A1(_10402_ ), .A2(_11278_ ), .A3(_11279_ ), .A4(_11296_ ), .ZN(_11297_ ) );
OAI21_X1 _15306_ ( .A(\u_lsu.pmem[6822] ), .B1(_11285_ ), .B2(_11293_ ), .ZN(_11298_ ) );
AOI21_X1 _15307_ ( .A(fanout_net_23 ), .B1(_11297_ ), .B2(_11298_ ), .ZN(_00628_ ) );
NAND4_X1 _15308_ ( .A1(_10405_ ), .A2(_11278_ ), .A3(_11279_ ), .A4(_11296_ ), .ZN(_11299_ ) );
OAI21_X1 _15309_ ( .A(\u_lsu.pmem[6821] ), .B1(_11285_ ), .B2(_11293_ ), .ZN(_11300_ ) );
AOI21_X1 _15310_ ( .A(fanout_net_23 ), .B1(_11299_ ), .B2(_11300_ ), .ZN(_00629_ ) );
BUF_X4 _15311_ ( .A(_10886_ ), .Z(_11301_ ) );
NAND4_X1 _15312_ ( .A1(_10339_ ), .A2(_11301_ ), .A3(_11279_ ), .A4(_11074_ ), .ZN(_11302_ ) );
OAI21_X1 _15313_ ( .A(\u_lsu.pmem[3812] ), .B1(_11214_ ), .B2(_10327_ ), .ZN(_11303_ ) );
AOI21_X1 _15314_ ( .A(fanout_net_23 ), .B1(_11302_ ), .B2(_11303_ ), .ZN(_00630_ ) );
NAND4_X1 _15315_ ( .A1(_10408_ ), .A2(_11278_ ), .A3(_11279_ ), .A4(_11296_ ), .ZN(_11304_ ) );
OAI21_X1 _15316_ ( .A(\u_lsu.pmem[6820] ), .B1(_11285_ ), .B2(_11293_ ), .ZN(_11305_ ) );
AOI21_X1 _15317_ ( .A(fanout_net_23 ), .B1(_11304_ ), .B2(_11305_ ), .ZN(_00631_ ) );
BUF_X4 _15318_ ( .A(_11063_ ), .Z(_11306_ ) );
NAND4_X1 _15319_ ( .A1(_10411_ ), .A2(_11278_ ), .A3(_11306_ ), .A4(_11296_ ), .ZN(_11307_ ) );
OAI21_X1 _15320_ ( .A(\u_lsu.pmem[6819] ), .B1(_11285_ ), .B2(_11293_ ), .ZN(_11308_ ) );
AOI21_X1 _15321_ ( .A(fanout_net_23 ), .B1(_11307_ ), .B2(_11308_ ), .ZN(_00632_ ) );
BUF_X4 _15322_ ( .A(_09671_ ), .Z(_11309_ ) );
NAND4_X1 _15323_ ( .A1(_10414_ ), .A2(_11309_ ), .A3(_11306_ ), .A4(_11296_ ), .ZN(_11310_ ) );
OAI21_X1 _15324_ ( .A(\u_lsu.pmem[6818] ), .B1(_11285_ ), .B2(_11293_ ), .ZN(_11311_ ) );
AOI21_X1 _15325_ ( .A(fanout_net_23 ), .B1(_11310_ ), .B2(_11311_ ), .ZN(_00633_ ) );
NAND4_X1 _15326_ ( .A1(_10417_ ), .A2(_11309_ ), .A3(_11306_ ), .A4(_11296_ ), .ZN(_11312_ ) );
OAI21_X1 _15327_ ( .A(\u_lsu.pmem[6817] ), .B1(_11285_ ), .B2(_11293_ ), .ZN(_11313_ ) );
AOI21_X1 _15328_ ( .A(fanout_net_23 ), .B1(_11312_ ), .B2(_11313_ ), .ZN(_00634_ ) );
OAI21_X1 _15329_ ( .A(\u_lsu.pmem[6816] ), .B1(_11218_ ), .B2(_11294_ ), .ZN(_11314_ ) );
NAND4_X1 _15330_ ( .A1(_10525_ ), .A2(_11061_ ), .A3(_11125_ ), .A4(_11292_ ), .ZN(_11315_ ) );
AOI21_X1 _15331_ ( .A(fanout_net_23 ), .B1(_11314_ ), .B2(_11315_ ), .ZN(_00635_ ) );
NAND3_X1 _15332_ ( .A1(_10423_ ), .A2(_09842_ ), .A3(_10424_ ), .ZN(_11316_ ) );
BUF_X4 _15333_ ( .A(_11316_ ), .Z(_11317_ ) );
OAI21_X1 _15334_ ( .A(\u_lsu.pmem[6791] ), .B1(_11317_ ), .B2(_11123_ ), .ZN(_11318_ ) );
NAND4_X1 _15335_ ( .A1(_10436_ ), .A2(_09540_ ), .A3(_11125_ ), .A4(_11128_ ), .ZN(_11319_ ) );
AOI21_X1 _15336_ ( .A(fanout_net_23 ), .B1(_11318_ ), .B2(_11319_ ), .ZN(_00636_ ) );
AND2_X2 _15337_ ( .A1(_10423_ ), .A2(_09539_ ), .ZN(_11320_ ) );
BUF_X4 _15338_ ( .A(_11320_ ), .Z(_11321_ ) );
NAND4_X1 _15339_ ( .A1(_11321_ ), .A2(_10444_ ), .A3(_11306_ ), .A4(_11296_ ), .ZN(_11322_ ) );
OAI21_X1 _15340_ ( .A(\u_lsu.pmem[6790] ), .B1(_11317_ ), .B2(_10465_ ), .ZN(_11323_ ) );
AOI21_X1 _15341_ ( .A(fanout_net_23 ), .B1(_11322_ ), .B2(_11323_ ), .ZN(_00637_ ) );
NAND4_X1 _15342_ ( .A1(_11321_ ), .A2(_10448_ ), .A3(_11306_ ), .A4(_11296_ ), .ZN(_11324_ ) );
OAI21_X1 _15343_ ( .A(\u_lsu.pmem[6789] ), .B1(_11317_ ), .B2(_10465_ ), .ZN(_11325_ ) );
AOI21_X1 _15344_ ( .A(fanout_net_24 ), .B1(_11324_ ), .B2(_11325_ ), .ZN(_00638_ ) );
NAND4_X1 _15345_ ( .A1(_11321_ ), .A2(_10453_ ), .A3(_11306_ ), .A4(_11296_ ), .ZN(_11326_ ) );
OAI21_X1 _15346_ ( .A(\u_lsu.pmem[6788] ), .B1(_11317_ ), .B2(_10465_ ), .ZN(_11327_ ) );
AOI21_X1 _15347_ ( .A(fanout_net_24 ), .B1(_11326_ ), .B2(_11327_ ), .ZN(_00639_ ) );
NAND4_X1 _15348_ ( .A1(_11321_ ), .A2(_10456_ ), .A3(_11306_ ), .A4(_11296_ ), .ZN(_11328_ ) );
OAI21_X1 _15349_ ( .A(\u_lsu.pmem[6787] ), .B1(_11317_ ), .B2(_10465_ ), .ZN(_11329_ ) );
AOI21_X1 _15350_ ( .A(fanout_net_24 ), .B1(_11328_ ), .B2(_11329_ ), .ZN(_00640_ ) );
NAND4_X1 _15351_ ( .A1(_10345_ ), .A2(_11301_ ), .A3(_11306_ ), .A4(_11074_ ), .ZN(_11330_ ) );
OAI21_X1 _15352_ ( .A(\u_lsu.pmem[3811] ), .B1(_11214_ ), .B2(_10327_ ), .ZN(_11331_ ) );
AOI21_X1 _15353_ ( .A(fanout_net_24 ), .B1(_11330_ ), .B2(_11331_ ), .ZN(_00641_ ) );
OAI21_X1 _15354_ ( .A(\u_lsu.pmem[6786] ), .B1(_11317_ ), .B2(_11123_ ), .ZN(_11332_ ) );
NAND4_X1 _15355_ ( .A1(_10460_ ), .A2(_09540_ ), .A3(_11125_ ), .A4(_11128_ ), .ZN(_11333_ ) );
AOI21_X1 _15356_ ( .A(fanout_net_24 ), .B1(_11332_ ), .B2(_11333_ ), .ZN(_00642_ ) );
BUF_X8 _15357_ ( .A(_09471_ ), .Z(_11334_ ) );
BUF_X4 _15358_ ( .A(_11334_ ), .Z(_11335_ ) );
NAND4_X1 _15359_ ( .A1(_11321_ ), .A2(_10463_ ), .A3(_11306_ ), .A4(_11335_ ), .ZN(_11336_ ) );
BUF_X4 _15360_ ( .A(_09515_ ), .Z(_11337_ ) );
OAI21_X1 _15361_ ( .A(\u_lsu.pmem[6785] ), .B1(_11317_ ), .B2(_11337_ ), .ZN(_11338_ ) );
AOI21_X1 _15362_ ( .A(fanout_net_24 ), .B1(_11336_ ), .B2(_11338_ ), .ZN(_00643_ ) );
NAND4_X1 _15363_ ( .A1(_11321_ ), .A2(_10467_ ), .A3(_11306_ ), .A4(_11335_ ), .ZN(_11339_ ) );
OAI21_X1 _15364_ ( .A(\u_lsu.pmem[6784] ), .B1(_11317_ ), .B2(_11337_ ), .ZN(_11340_ ) );
AOI21_X1 _15365_ ( .A(fanout_net_24 ), .B1(_11339_ ), .B2(_11340_ ), .ZN(_00644_ ) );
NOR2_X2 _15366_ ( .A1(_10470_ ), .A2(_09118_ ), .ZN(_11341_ ) );
NAND2_X1 _15367_ ( .A1(_11341_ ), .A2(_10325_ ), .ZN(_11342_ ) );
BUF_X4 _15368_ ( .A(_11342_ ), .Z(_11343_ ) );
OAI21_X1 _15369_ ( .A(\u_lsu.pmem[6759] ), .B1(_11218_ ), .B2(_11343_ ), .ZN(_11344_ ) );
NAND4_X1 _15370_ ( .A1(_10851_ ), .A2(_11061_ ), .A3(_11125_ ), .A4(_11341_ ), .ZN(_11345_ ) );
AOI21_X1 _15371_ ( .A(fanout_net_24 ), .B1(_11344_ ), .B2(_11345_ ), .ZN(_00645_ ) );
OAI21_X1 _15372_ ( .A(\u_lsu.pmem[6758] ), .B1(_11218_ ), .B2(_11343_ ), .ZN(_11346_ ) );
BUF_X4 _15373_ ( .A(_09578_ ), .Z(_11347_ ) );
BUF_X4 _15374_ ( .A(_09878_ ), .Z(_11348_ ) );
NAND4_X1 _15375_ ( .A1(_11347_ ), .A2(_11061_ ), .A3(_11348_ ), .A4(_11341_ ), .ZN(_11349_ ) );
AOI21_X1 _15376_ ( .A(fanout_net_24 ), .B1(_11346_ ), .B2(_11349_ ), .ZN(_00646_ ) );
OAI21_X1 _15377_ ( .A(\u_lsu.pmem[6757] ), .B1(_11218_ ), .B2(_11343_ ), .ZN(_11350_ ) );
BUF_X4 _15378_ ( .A(_09585_ ), .Z(_11351_ ) );
NAND4_X1 _15379_ ( .A1(_11351_ ), .A2(_11061_ ), .A3(_11348_ ), .A4(_11341_ ), .ZN(_11352_ ) );
AOI21_X1 _15380_ ( .A(fanout_net_24 ), .B1(_11350_ ), .B2(_11352_ ), .ZN(_00647_ ) );
OAI21_X1 _15381_ ( .A(\u_lsu.pmem[6756] ), .B1(_11218_ ), .B2(_11343_ ), .ZN(_11353_ ) );
NAND4_X1 _15382_ ( .A1(_10486_ ), .A2(_11061_ ), .A3(_11348_ ), .A4(_11341_ ), .ZN(_11354_ ) );
AOI21_X1 _15383_ ( .A(fanout_net_24 ), .B1(_11353_ ), .B2(_11354_ ), .ZN(_00648_ ) );
OAI21_X1 _15384_ ( .A(\u_lsu.pmem[6755] ), .B1(_11218_ ), .B2(_11343_ ), .ZN(_11355_ ) );
NAND4_X1 _15385_ ( .A1(_09449_ ), .A2(_11061_ ), .A3(_11348_ ), .A4(_11341_ ), .ZN(_11356_ ) );
AOI21_X1 _15386_ ( .A(fanout_net_24 ), .B1(_11355_ ), .B2(_11356_ ), .ZN(_00649_ ) );
BUF_X4 _15387_ ( .A(_09572_ ), .Z(_11357_ ) );
OAI21_X1 _15388_ ( .A(\u_lsu.pmem[6754] ), .B1(_11357_ ), .B2(_11343_ ), .ZN(_11358_ ) );
BUF_X4 _15389_ ( .A(_10548_ ), .Z(_11359_ ) );
NAND4_X1 _15390_ ( .A1(_10492_ ), .A2(_11359_ ), .A3(_11348_ ), .A4(_11341_ ), .ZN(_11360_ ) );
AOI21_X1 _15391_ ( .A(fanout_net_24 ), .B1(_11358_ ), .B2(_11360_ ), .ZN(_00650_ ) );
OAI21_X1 _15392_ ( .A(\u_lsu.pmem[6753] ), .B1(_11357_ ), .B2(_11343_ ), .ZN(_11361_ ) );
NAND4_X1 _15393_ ( .A1(_09698_ ), .A2(_11359_ ), .A3(_11348_ ), .A4(_11341_ ), .ZN(_11362_ ) );
AOI21_X1 _15394_ ( .A(fanout_net_24 ), .B1(_11361_ ), .B2(_11362_ ), .ZN(_00651_ ) );
BUF_X4 _15395_ ( .A(_11063_ ), .Z(_11363_ ) );
NAND4_X1 _15396_ ( .A1(_10350_ ), .A2(_11301_ ), .A3(_11363_ ), .A4(_11074_ ), .ZN(_11364_ ) );
OAI21_X1 _15397_ ( .A(\u_lsu.pmem[3810] ), .B1(_11214_ ), .B2(_10327_ ), .ZN(_11365_ ) );
AOI21_X1 _15398_ ( .A(fanout_net_24 ), .B1(_11364_ ), .B2(_11365_ ), .ZN(_00652_ ) );
OAI21_X1 _15399_ ( .A(\u_lsu.pmem[6752] ), .B1(_11357_ ), .B2(_11343_ ), .ZN(_11366_ ) );
NAND4_X1 _15400_ ( .A1(_10525_ ), .A2(_11359_ ), .A3(_11348_ ), .A4(_11341_ ), .ZN(_11367_ ) );
AOI21_X1 _15401_ ( .A(fanout_net_24 ), .B1(_11366_ ), .B2(_11367_ ), .ZN(_00653_ ) );
AND3_X1 _15402_ ( .A1(_09506_ ), .A2(_09130_ ), .A3(_09947_ ), .ZN(_11368_ ) );
BUF_X4 _15403_ ( .A(_11368_ ), .Z(_11369_ ) );
NAND2_X1 _15404_ ( .A1(_11369_ ), .A2(_11028_ ), .ZN(_11370_ ) );
BUF_X4 _15405_ ( .A(_11370_ ), .Z(_11371_ ) );
OAI21_X1 _15406_ ( .A(\u_lsu.pmem[6727] ), .B1(_11357_ ), .B2(_11371_ ), .ZN(_11372_ ) );
BUF_X4 _15407_ ( .A(_11369_ ), .Z(_11373_ ) );
NAND4_X1 _15408_ ( .A1(_10851_ ), .A2(_11359_ ), .A3(_11348_ ), .A4(_11373_ ), .ZN(_11374_ ) );
AOI21_X1 _15409_ ( .A(fanout_net_24 ), .B1(_11372_ ), .B2(_11374_ ), .ZN(_00654_ ) );
OAI21_X1 _15410_ ( .A(\u_lsu.pmem[6726] ), .B1(_11357_ ), .B2(_11371_ ), .ZN(_11375_ ) );
NAND4_X1 _15411_ ( .A1(_11347_ ), .A2(_11359_ ), .A3(_11348_ ), .A4(_11373_ ), .ZN(_11376_ ) );
AOI21_X1 _15412_ ( .A(fanout_net_24 ), .B1(_11375_ ), .B2(_11376_ ), .ZN(_00655_ ) );
OAI21_X1 _15413_ ( .A(\u_lsu.pmem[6725] ), .B1(_11357_ ), .B2(_11370_ ), .ZN(_11377_ ) );
BUF_X4 _15414_ ( .A(_11369_ ), .Z(_11378_ ) );
NAND4_X1 _15415_ ( .A1(_11351_ ), .A2(_11359_ ), .A3(_11348_ ), .A4(_11378_ ), .ZN(_11379_ ) );
AOI21_X1 _15416_ ( .A(fanout_net_24 ), .B1(_11377_ ), .B2(_11379_ ), .ZN(_00656_ ) );
OAI21_X1 _15417_ ( .A(\u_lsu.pmem[6724] ), .B1(_11357_ ), .B2(_11370_ ), .ZN(_11380_ ) );
BUF_X8 _15418_ ( .A(_09877_ ), .Z(_11381_ ) );
BUF_X4 _15419_ ( .A(_11381_ ), .Z(_11382_ ) );
NAND4_X1 _15420_ ( .A1(_10486_ ), .A2(_11359_ ), .A3(_11382_ ), .A4(_11378_ ), .ZN(_11383_ ) );
AOI21_X1 _15421_ ( .A(fanout_net_24 ), .B1(_11380_ ), .B2(_11383_ ), .ZN(_00657_ ) );
OAI21_X1 _15422_ ( .A(\u_lsu.pmem[6723] ), .B1(_11357_ ), .B2(_11370_ ), .ZN(_11384_ ) );
BUF_X4 _15423_ ( .A(_09448_ ), .Z(_11385_ ) );
NAND4_X1 _15424_ ( .A1(_11385_ ), .A2(_11359_ ), .A3(_11382_ ), .A4(_11378_ ), .ZN(_11386_ ) );
AOI21_X1 _15425_ ( .A(fanout_net_24 ), .B1(_11384_ ), .B2(_11386_ ), .ZN(_00658_ ) );
OAI21_X1 _15426_ ( .A(\u_lsu.pmem[6722] ), .B1(_11357_ ), .B2(_11370_ ), .ZN(_11387_ ) );
NAND4_X1 _15427_ ( .A1(_10492_ ), .A2(_11359_ ), .A3(_11382_ ), .A4(_11378_ ), .ZN(_11388_ ) );
AOI21_X1 _15428_ ( .A(fanout_net_24 ), .B1(_11387_ ), .B2(_11388_ ), .ZN(_00659_ ) );
OAI21_X1 _15429_ ( .A(\u_lsu.pmem[6721] ), .B1(_11357_ ), .B2(_11370_ ), .ZN(_11389_ ) );
NAND4_X1 _15430_ ( .A1(_09698_ ), .A2(_11359_ ), .A3(_11382_ ), .A4(_11378_ ), .ZN(_11390_ ) );
AOI21_X1 _15431_ ( .A(fanout_net_24 ), .B1(_11389_ ), .B2(_11390_ ), .ZN(_00660_ ) );
BUF_X4 _15432_ ( .A(_09572_ ), .Z(_11391_ ) );
OAI21_X1 _15433_ ( .A(\u_lsu.pmem[6720] ), .B1(_11391_ ), .B2(_11370_ ), .ZN(_11392_ ) );
BUF_X4 _15434_ ( .A(_10548_ ), .Z(_11393_ ) );
NAND4_X1 _15435_ ( .A1(_10525_ ), .A2(_11393_ ), .A3(_11382_ ), .A4(_11378_ ), .ZN(_11394_ ) );
AOI21_X1 _15436_ ( .A(fanout_net_24 ), .B1(_11392_ ), .B2(_11394_ ), .ZN(_00661_ ) );
NAND4_X1 _15437_ ( .A1(_10527_ ), .A2(_11309_ ), .A3(_11363_ ), .A4(_11335_ ), .ZN(_11395_ ) );
BUF_X4 _15438_ ( .A(_10844_ ), .Z(_11396_ ) );
NAND3_X1 _15439_ ( .A1(_09135_ ), .A2(_09538_ ), .A3(_10530_ ), .ZN(_11397_ ) );
BUF_X4 _15440_ ( .A(_11397_ ), .Z(_11398_ ) );
OAI21_X1 _15441_ ( .A(\u_lsu.pmem[6695] ), .B1(_11396_ ), .B2(_11398_ ), .ZN(_11399_ ) );
AOI21_X1 _15442_ ( .A(fanout_net_24 ), .B1(_11395_ ), .B2(_11399_ ), .ZN(_00662_ ) );
NAND4_X1 _15443_ ( .A1(_10354_ ), .A2(_11301_ ), .A3(_11363_ ), .A4(_11074_ ), .ZN(_11400_ ) );
OAI21_X1 _15444_ ( .A(\u_lsu.pmem[3809] ), .B1(_11214_ ), .B2(_10327_ ), .ZN(_11401_ ) );
AOI21_X1 _15445_ ( .A(fanout_net_24 ), .B1(_11400_ ), .B2(_11401_ ), .ZN(_00663_ ) );
NAND4_X1 _15446_ ( .A1(_10535_ ), .A2(_11309_ ), .A3(_11363_ ), .A4(_11335_ ), .ZN(_11402_ ) );
OAI21_X1 _15447_ ( .A(\u_lsu.pmem[6694] ), .B1(_11396_ ), .B2(_11398_ ), .ZN(_11403_ ) );
AOI21_X1 _15448_ ( .A(fanout_net_24 ), .B1(_11402_ ), .B2(_11403_ ), .ZN(_00664_ ) );
NAND4_X1 _15449_ ( .A1(_10538_ ), .A2(_11309_ ), .A3(_11363_ ), .A4(_11335_ ), .ZN(_11404_ ) );
OAI21_X1 _15450_ ( .A(\u_lsu.pmem[6693] ), .B1(_11396_ ), .B2(_11398_ ), .ZN(_11405_ ) );
AOI21_X1 _15451_ ( .A(fanout_net_24 ), .B1(_11404_ ), .B2(_11405_ ), .ZN(_00665_ ) );
OAI21_X1 _15452_ ( .A(\u_lsu.pmem[6692] ), .B1(_11391_ ), .B2(_11398_ ), .ZN(_11406_ ) );
AND2_X1 _15453_ ( .A1(_09539_ ), .A2(_10530_ ), .ZN(_11407_ ) );
NAND4_X1 _15454_ ( .A1(_10486_ ), .A2(_11393_ ), .A3(_11382_ ), .A4(_11407_ ), .ZN(_11408_ ) );
AOI21_X1 _15455_ ( .A(fanout_net_24 ), .B1(_11406_ ), .B2(_11408_ ), .ZN(_00666_ ) );
OAI21_X1 _15456_ ( .A(\u_lsu.pmem[6691] ), .B1(_11391_ ), .B2(_11398_ ), .ZN(_11409_ ) );
NAND4_X1 _15457_ ( .A1(_11385_ ), .A2(_11393_ ), .A3(_11382_ ), .A4(_11407_ ), .ZN(_11410_ ) );
AOI21_X1 _15458_ ( .A(fanout_net_24 ), .B1(_11409_ ), .B2(_11410_ ), .ZN(_00667_ ) );
OAI21_X1 _15459_ ( .A(\u_lsu.pmem[6690] ), .B1(_11391_ ), .B2(_11398_ ), .ZN(_11411_ ) );
NAND4_X1 _15460_ ( .A1(_10492_ ), .A2(_11393_ ), .A3(_11382_ ), .A4(_11407_ ), .ZN(_11412_ ) );
AOI21_X1 _15461_ ( .A(fanout_net_25 ), .B1(_11411_ ), .B2(_11412_ ), .ZN(_00668_ ) );
OAI21_X1 _15462_ ( .A(\u_lsu.pmem[6689] ), .B1(_11391_ ), .B2(_11398_ ), .ZN(_11413_ ) );
BUF_X4 _15463_ ( .A(_09616_ ), .Z(_11414_ ) );
NAND4_X1 _15464_ ( .A1(_11414_ ), .A2(_11393_ ), .A3(_11382_ ), .A4(_11407_ ), .ZN(_11415_ ) );
AOI21_X1 _15465_ ( .A(fanout_net_25 ), .B1(_11413_ ), .B2(_11415_ ), .ZN(_00669_ ) );
NAND4_X1 _15466_ ( .A1(_10556_ ), .A2(_11309_ ), .A3(_11363_ ), .A4(_11335_ ), .ZN(_11416_ ) );
OAI21_X1 _15467_ ( .A(\u_lsu.pmem[6688] ), .B1(_11396_ ), .B2(_11398_ ), .ZN(_11417_ ) );
AOI21_X1 _15468_ ( .A(fanout_net_25 ), .B1(_11416_ ), .B2(_11417_ ), .ZN(_00670_ ) );
AND3_X1 _15469_ ( .A1(_09135_ ), .A2(_10560_ ), .A3(_09538_ ), .ZN(_11418_ ) );
INV_X1 _15470_ ( .A(_11418_ ), .ZN(_11419_ ) );
BUF_X4 _15471_ ( .A(_11419_ ), .Z(_11420_ ) );
OAI21_X1 _15472_ ( .A(\u_lsu.pmem[6663] ), .B1(_11420_ ), .B2(_11123_ ), .ZN(_11421_ ) );
BUF_X4 _15473_ ( .A(_11418_ ), .Z(_11422_ ) );
BUF_X4 _15474_ ( .A(_08582_ ), .Z(_11423_ ) );
NAND3_X1 _15475_ ( .A1(_11422_ ), .A2(_11423_ ), .A3(_10785_ ), .ZN(_11424_ ) );
AOI21_X1 _15476_ ( .A(fanout_net_25 ), .B1(_11421_ ), .B2(_11424_ ), .ZN(_00671_ ) );
OAI21_X1 _15477_ ( .A(\u_lsu.pmem[6662] ), .B1(_11420_ ), .B2(_11123_ ), .ZN(_11425_ ) );
BUF_X4 _15478_ ( .A(_09472_ ), .Z(_11426_ ) );
NAND3_X1 _15479_ ( .A1(_11422_ ), .A2(_10444_ ), .A3(_11426_ ), .ZN(_11427_ ) );
AOI21_X1 _15480_ ( .A(fanout_net_25 ), .B1(_11425_ ), .B2(_11427_ ), .ZN(_00672_ ) );
OAI21_X1 _15481_ ( .A(\u_lsu.pmem[6661] ), .B1(_11420_ ), .B2(_11123_ ), .ZN(_11428_ ) );
NAND3_X1 _15482_ ( .A1(_11422_ ), .A2(_10448_ ), .A3(_11426_ ), .ZN(_11429_ ) );
AOI21_X1 _15483_ ( .A(fanout_net_25 ), .B1(_11428_ ), .B2(_11429_ ), .ZN(_00673_ ) );
NAND4_X1 _15484_ ( .A1(_10357_ ), .A2(_11301_ ), .A3(_11363_ ), .A4(_11074_ ), .ZN(_11430_ ) );
OAI21_X1 _15485_ ( .A(\u_lsu.pmem[3808] ), .B1(_11214_ ), .B2(_10327_ ), .ZN(_11431_ ) );
AOI21_X1 _15486_ ( .A(fanout_net_25 ), .B1(_11430_ ), .B2(_11431_ ), .ZN(_00674_ ) );
OAI21_X1 _15487_ ( .A(\u_lsu.pmem[6660] ), .B1(_11420_ ), .B2(_11123_ ), .ZN(_11432_ ) );
NAND3_X1 _15488_ ( .A1(_11422_ ), .A2(_10453_ ), .A3(_11426_ ), .ZN(_11433_ ) );
AOI21_X1 _15489_ ( .A(fanout_net_25 ), .B1(_11432_ ), .B2(_11433_ ), .ZN(_00675_ ) );
NAND4_X1 _15490_ ( .A1(_10575_ ), .A2(_11309_ ), .A3(_11363_ ), .A4(_11335_ ), .ZN(_11434_ ) );
OAI21_X1 _15491_ ( .A(\u_lsu.pmem[6659] ), .B1(_11419_ ), .B2(_11337_ ), .ZN(_11435_ ) );
AOI21_X1 _15492_ ( .A(fanout_net_25 ), .B1(_11434_ ), .B2(_11435_ ), .ZN(_00676_ ) );
NAND4_X1 _15493_ ( .A1(_10584_ ), .A2(_09806_ ), .A3(_11363_ ), .A4(_11335_ ), .ZN(_11436_ ) );
OAI21_X1 _15494_ ( .A(\u_lsu.pmem[6658] ), .B1(_11419_ ), .B2(_11337_ ), .ZN(_11437_ ) );
AOI21_X1 _15495_ ( .A(fanout_net_25 ), .B1(_11436_ ), .B2(_11437_ ), .ZN(_00677_ ) );
OAI21_X1 _15496_ ( .A(\u_lsu.pmem[6657] ), .B1(_11420_ ), .B2(_11123_ ), .ZN(_11438_ ) );
NAND3_X1 _15497_ ( .A1(_11422_ ), .A2(_10463_ ), .A3(_11426_ ), .ZN(_11439_ ) );
AOI21_X1 _15498_ ( .A(fanout_net_25 ), .B1(_11438_ ), .B2(_11439_ ), .ZN(_00678_ ) );
NAND4_X1 _15499_ ( .A1(_10591_ ), .A2(_11309_ ), .A3(_11363_ ), .A4(_11335_ ), .ZN(_11440_ ) );
OAI21_X1 _15500_ ( .A(\u_lsu.pmem[6656] ), .B1(_11419_ ), .B2(_11337_ ), .ZN(_11441_ ) );
AOI21_X1 _15501_ ( .A(fanout_net_25 ), .B1(_11440_ ), .B2(_11441_ ), .ZN(_00679_ ) );
NOR3_X4 _15502_ ( .A1(_10397_ ), .A2(_09462_ ), .A3(_11029_ ), .ZN(_11442_ ) );
NAND2_X2 _15503_ ( .A1(_11442_ ), .A2(_10424_ ), .ZN(_11443_ ) );
BUF_X4 _15504_ ( .A(_11443_ ), .Z(_11444_ ) );
OAI21_X1 _15505_ ( .A(\u_lsu.pmem[6631] ), .B1(_11391_ ), .B2(_11444_ ), .ZN(_11445_ ) );
NAND4_X1 _15506_ ( .A1(_10851_ ), .A2(_11393_ ), .A3(_11382_ ), .A4(_11442_ ), .ZN(_11446_ ) );
AOI21_X1 _15507_ ( .A(fanout_net_25 ), .B1(_11445_ ), .B2(_11446_ ), .ZN(_00680_ ) );
BUF_X4 _15508_ ( .A(_11063_ ), .Z(_11447_ ) );
NAND4_X1 _15509_ ( .A1(_10603_ ), .A2(_11309_ ), .A3(_11447_ ), .A4(_11335_ ), .ZN(_11448_ ) );
OAI21_X1 _15510_ ( .A(\u_lsu.pmem[6630] ), .B1(_11396_ ), .B2(_11444_ ), .ZN(_11449_ ) );
AOI21_X1 _15511_ ( .A(fanout_net_25 ), .B1(_11448_ ), .B2(_11449_ ), .ZN(_00681_ ) );
BUF_X4 _15512_ ( .A(_11334_ ), .Z(_11450_ ) );
NAND4_X1 _15513_ ( .A1(_10608_ ), .A2(_11309_ ), .A3(_11447_ ), .A4(_11450_ ), .ZN(_11451_ ) );
OAI21_X1 _15514_ ( .A(\u_lsu.pmem[6629] ), .B1(_11396_ ), .B2(_11444_ ), .ZN(_11452_ ) );
AOI21_X1 _15515_ ( .A(fanout_net_25 ), .B1(_11451_ ), .B2(_11452_ ), .ZN(_00682_ ) );
BUF_X8 _15516_ ( .A(_09539_ ), .Z(_11453_ ) );
BUF_X4 _15517_ ( .A(_11453_ ), .Z(_11454_ ) );
NAND4_X1 _15518_ ( .A1(_10611_ ), .A2(_11454_ ), .A3(_11447_ ), .A4(_11450_ ), .ZN(_11455_ ) );
OAI21_X1 _15519_ ( .A(\u_lsu.pmem[6628] ), .B1(_11396_ ), .B2(_11444_ ), .ZN(_11456_ ) );
AOI21_X1 _15520_ ( .A(fanout_net_25 ), .B1(_11455_ ), .B2(_11456_ ), .ZN(_00683_ ) );
NAND4_X1 _15521_ ( .A1(_10614_ ), .A2(_11454_ ), .A3(_11447_ ), .A4(_11450_ ), .ZN(_11457_ ) );
OAI21_X1 _15522_ ( .A(\u_lsu.pmem[6627] ), .B1(_11396_ ), .B2(_11444_ ), .ZN(_11458_ ) );
AOI21_X1 _15523_ ( .A(fanout_net_25 ), .B1(_11457_ ), .B2(_11458_ ), .ZN(_00684_ ) );
NAND4_X1 _15524_ ( .A1(_10018_ ), .A2(_11212_ ), .A3(_09914_ ), .A4(_10362_ ), .ZN(_11459_ ) );
BUF_X4 _15525_ ( .A(_09562_ ), .Z(_11460_ ) );
OAI21_X1 _15526_ ( .A(\u_lsu.pmem[3783] ), .B1(_11460_ ), .B2(_10364_ ), .ZN(_11461_ ) );
AOI21_X1 _15527_ ( .A(fanout_net_25 ), .B1(_11459_ ), .B2(_11461_ ), .ZN(_00685_ ) );
NAND4_X1 _15528_ ( .A1(_10617_ ), .A2(_11454_ ), .A3(_11447_ ), .A4(_11450_ ), .ZN(_11462_ ) );
OAI21_X1 _15529_ ( .A(\u_lsu.pmem[6626] ), .B1(_11396_ ), .B2(_11444_ ), .ZN(_11463_ ) );
AOI21_X1 _15530_ ( .A(fanout_net_25 ), .B1(_11462_ ), .B2(_11463_ ), .ZN(_00686_ ) );
NAND4_X1 _15531_ ( .A1(_10621_ ), .A2(_11454_ ), .A3(_11447_ ), .A4(_11450_ ), .ZN(_11464_ ) );
OAI21_X1 _15532_ ( .A(\u_lsu.pmem[6625] ), .B1(_11396_ ), .B2(_11444_ ), .ZN(_11465_ ) );
AOI21_X1 _15533_ ( .A(fanout_net_25 ), .B1(_11464_ ), .B2(_11465_ ), .ZN(_00687_ ) );
NAND4_X1 _15534_ ( .A1(_10624_ ), .A2(_11454_ ), .A3(_11447_ ), .A4(_11450_ ), .ZN(_11466_ ) );
BUF_X4 _15535_ ( .A(_10844_ ), .Z(_11467_ ) );
OAI21_X1 _15536_ ( .A(\u_lsu.pmem[6624] ), .B1(_11467_ ), .B2(_11444_ ), .ZN(_11468_ ) );
AOI21_X1 _15537_ ( .A(fanout_net_25 ), .B1(_11466_ ), .B2(_11468_ ), .ZN(_00688_ ) );
NOR3_X4 _15538_ ( .A1(_10397_ ), .A2(_09462_ ), .A3(_11055_ ), .ZN(_11469_ ) );
NAND2_X2 _15539_ ( .A1(_11469_ ), .A2(_10424_ ), .ZN(_11470_ ) );
BUF_X4 _15540_ ( .A(_11470_ ), .Z(_11471_ ) );
OAI21_X1 _15541_ ( .A(\u_lsu.pmem[6599] ), .B1(_11391_ ), .B2(_11471_ ), .ZN(_11472_ ) );
BUF_X4 _15542_ ( .A(_11381_ ), .Z(_11473_ ) );
NAND4_X1 _15543_ ( .A1(_10851_ ), .A2(_11393_ ), .A3(_11473_ ), .A4(_11469_ ), .ZN(_11474_ ) );
AOI21_X1 _15544_ ( .A(fanout_net_25 ), .B1(_11472_ ), .B2(_11474_ ), .ZN(_00689_ ) );
NAND4_X1 _15545_ ( .A1(_10632_ ), .A2(_11454_ ), .A3(_11447_ ), .A4(_11450_ ), .ZN(_11475_ ) );
OAI21_X1 _15546_ ( .A(\u_lsu.pmem[6598] ), .B1(_11467_ ), .B2(_11471_ ), .ZN(_11476_ ) );
AOI21_X1 _15547_ ( .A(fanout_net_25 ), .B1(_11475_ ), .B2(_11476_ ), .ZN(_00690_ ) );
NAND4_X1 _15548_ ( .A1(_10635_ ), .A2(_11454_ ), .A3(_11447_ ), .A4(_11450_ ), .ZN(_11477_ ) );
OAI21_X1 _15549_ ( .A(\u_lsu.pmem[6597] ), .B1(_11467_ ), .B2(_11471_ ), .ZN(_11478_ ) );
AOI21_X1 _15550_ ( .A(fanout_net_25 ), .B1(_11477_ ), .B2(_11478_ ), .ZN(_00691_ ) );
NAND4_X1 _15551_ ( .A1(_10641_ ), .A2(_11454_ ), .A3(_11447_ ), .A4(_11450_ ), .ZN(_11479_ ) );
OAI21_X1 _15552_ ( .A(\u_lsu.pmem[6596] ), .B1(_11467_ ), .B2(_11471_ ), .ZN(_11480_ ) );
AOI21_X1 _15553_ ( .A(fanout_net_25 ), .B1(_11479_ ), .B2(_11480_ ), .ZN(_00692_ ) );
BUF_X4 _15554_ ( .A(_11063_ ), .Z(_11481_ ) );
NAND4_X1 _15555_ ( .A1(_10645_ ), .A2(_11454_ ), .A3(_11481_ ), .A4(_11450_ ), .ZN(_11482_ ) );
OAI21_X1 _15556_ ( .A(\u_lsu.pmem[6595] ), .B1(_11467_ ), .B2(_11471_ ), .ZN(_11483_ ) );
AOI21_X1 _15557_ ( .A(fanout_net_25 ), .B1(_11482_ ), .B2(_11483_ ), .ZN(_00693_ ) );
BUF_X4 _15558_ ( .A(_11334_ ), .Z(_11484_ ) );
NAND4_X1 _15559_ ( .A1(_10649_ ), .A2(_11454_ ), .A3(_11481_ ), .A4(_11484_ ), .ZN(_11485_ ) );
OAI21_X1 _15560_ ( .A(\u_lsu.pmem[6594] ), .B1(_11467_ ), .B2(_11471_ ), .ZN(_11486_ ) );
AOI21_X1 _15561_ ( .A(fanout_net_25 ), .B1(_11485_ ), .B2(_11486_ ), .ZN(_00694_ ) );
BUF_X4 _15562_ ( .A(_11453_ ), .Z(_11487_ ) );
NAND4_X1 _15563_ ( .A1(_10652_ ), .A2(_11487_ ), .A3(_11481_ ), .A4(_11484_ ), .ZN(_11488_ ) );
OAI21_X1 _15564_ ( .A(\u_lsu.pmem[6593] ), .B1(_11467_ ), .B2(_11471_ ), .ZN(_11489_ ) );
AOI21_X1 _15565_ ( .A(fanout_net_25 ), .B1(_11488_ ), .B2(_11489_ ), .ZN(_00695_ ) );
NAND4_X1 _15566_ ( .A1(_09763_ ), .A2(_11487_ ), .A3(_09869_ ), .A4(_11484_ ), .ZN(_11490_ ) );
OAI21_X1 _15567_ ( .A(\u_lsu.pmem[4325] ), .B1(_11467_ ), .B2(_09751_ ), .ZN(_11491_ ) );
AOI21_X1 _15568_ ( .A(fanout_net_25 ), .B1(_11490_ ), .B2(_11491_ ), .ZN(_00696_ ) );
BUF_X8 _15569_ ( .A(_09442_ ), .Z(_11492_ ) );
BUF_X4 _15570_ ( .A(_11492_ ), .Z(_11493_ ) );
NAND4_X1 _15571_ ( .A1(_10368_ ), .A2(_11301_ ), .A3(_11481_ ), .A4(_11493_ ), .ZN(_11494_ ) );
OAI21_X1 _15572_ ( .A(\u_lsu.pmem[3782] ), .B1(_11460_ ), .B2(_10364_ ), .ZN(_11495_ ) );
AOI21_X1 _15573_ ( .A(fanout_net_25 ), .B1(_11494_ ), .B2(_11495_ ), .ZN(_00697_ ) );
NAND4_X1 _15574_ ( .A1(_10655_ ), .A2(_11487_ ), .A3(_11481_ ), .A4(_11484_ ), .ZN(_11496_ ) );
OAI21_X1 _15575_ ( .A(\u_lsu.pmem[6592] ), .B1(_11467_ ), .B2(_11471_ ), .ZN(_11497_ ) );
AOI21_X1 _15576_ ( .A(fanout_net_26 ), .B1(_11496_ ), .B2(_11497_ ), .ZN(_00698_ ) );
NAND4_X1 _15577_ ( .A1(_10658_ ), .A2(_11487_ ), .A3(_11481_ ), .A4(_11484_ ), .ZN(_11498_ ) );
AND3_X2 _15578_ ( .A1(_09506_ ), .A2(_09505_ ), .A3(_10165_ ), .ZN(_11499_ ) );
NAND2_X1 _15579_ ( .A1(_11499_ ), .A2(_11028_ ), .ZN(_11500_ ) );
BUF_X4 _15580_ ( .A(_11500_ ), .Z(_11501_ ) );
OAI21_X1 _15581_ ( .A(\u_lsu.pmem[6567] ), .B1(_11467_ ), .B2(_11501_ ), .ZN(_11502_ ) );
AOI21_X1 _15582_ ( .A(fanout_net_26 ), .B1(_11498_ ), .B2(_11502_ ), .ZN(_00699_ ) );
NAND4_X1 _15583_ ( .A1(_10665_ ), .A2(_11487_ ), .A3(_11481_ ), .A4(_11484_ ), .ZN(_11503_ ) );
BUF_X4 _15584_ ( .A(_10844_ ), .Z(_11504_ ) );
OAI21_X1 _15585_ ( .A(\u_lsu.pmem[6566] ), .B1(_11504_ ), .B2(_11500_ ), .ZN(_11505_ ) );
AOI21_X1 _15586_ ( .A(fanout_net_26 ), .B1(_11503_ ), .B2(_11505_ ), .ZN(_00700_ ) );
NAND4_X1 _15587_ ( .A1(_10668_ ), .A2(_11487_ ), .A3(_11481_ ), .A4(_11484_ ), .ZN(_11506_ ) );
OAI21_X1 _15588_ ( .A(\u_lsu.pmem[6565] ), .B1(_11504_ ), .B2(_11500_ ), .ZN(_11507_ ) );
AOI21_X1 _15589_ ( .A(fanout_net_26 ), .B1(_11506_ ), .B2(_11507_ ), .ZN(_00701_ ) );
NAND4_X1 _15590_ ( .A1(_10671_ ), .A2(_11487_ ), .A3(_11481_ ), .A4(_11484_ ), .ZN(_11508_ ) );
OAI21_X1 _15591_ ( .A(\u_lsu.pmem[6564] ), .B1(_11504_ ), .B2(_11500_ ), .ZN(_11509_ ) );
AOI21_X1 _15592_ ( .A(fanout_net_26 ), .B1(_11508_ ), .B2(_11509_ ), .ZN(_00702_ ) );
NAND4_X1 _15593_ ( .A1(_10674_ ), .A2(_11487_ ), .A3(_11481_ ), .A4(_11484_ ), .ZN(_11510_ ) );
OAI21_X1 _15594_ ( .A(\u_lsu.pmem[6563] ), .B1(_11504_ ), .B2(_11500_ ), .ZN(_11511_ ) );
AOI21_X1 _15595_ ( .A(fanout_net_26 ), .B1(_11510_ ), .B2(_11511_ ), .ZN(_00703_ ) );
BUF_X4 _15596_ ( .A(_11063_ ), .Z(_11512_ ) );
NAND4_X1 _15597_ ( .A1(_10679_ ), .A2(_11487_ ), .A3(_11512_ ), .A4(_11484_ ), .ZN(_11513_ ) );
OAI21_X1 _15598_ ( .A(\u_lsu.pmem[6562] ), .B1(_11504_ ), .B2(_11500_ ), .ZN(_11514_ ) );
AOI21_X1 _15599_ ( .A(fanout_net_26 ), .B1(_11513_ ), .B2(_11514_ ), .ZN(_00704_ ) );
BUF_X4 _15600_ ( .A(_11334_ ), .Z(_11515_ ) );
NAND4_X1 _15601_ ( .A1(_10682_ ), .A2(_11487_ ), .A3(_11512_ ), .A4(_11515_ ), .ZN(_11516_ ) );
OAI21_X1 _15602_ ( .A(\u_lsu.pmem[6561] ), .B1(_11504_ ), .B2(_11500_ ), .ZN(_11517_ ) );
AOI21_X1 _15603_ ( .A(fanout_net_26 ), .B1(_11516_ ), .B2(_11517_ ), .ZN(_00705_ ) );
OAI21_X1 _15604_ ( .A(\u_lsu.pmem[6560] ), .B1(_11391_ ), .B2(_11501_ ), .ZN(_11518_ ) );
NAND4_X1 _15605_ ( .A1(_10525_ ), .A2(_11393_ ), .A3(_11473_ ), .A4(_11499_ ), .ZN(_11519_ ) );
AOI21_X1 _15606_ ( .A(fanout_net_26 ), .B1(_11518_ ), .B2(_11519_ ), .ZN(_00706_ ) );
NAND2_X1 _15607_ ( .A1(_09507_ ), .A2(_11028_ ), .ZN(_11520_ ) );
BUF_X4 _15608_ ( .A(_11520_ ), .Z(_11521_ ) );
BUF_X4 _15609_ ( .A(_10901_ ), .Z(_11522_ ) );
OAI21_X1 _15610_ ( .A(\u_lsu.pmem[6535] ), .B1(_11521_ ), .B2(_11522_ ), .ZN(_11523_ ) );
NAND4_X1 _15611_ ( .A1(_09513_ ), .A2(_10752_ ), .A3(_11473_ ), .A4(_11128_ ), .ZN(_11524_ ) );
AOI21_X1 _15612_ ( .A(fanout_net_26 ), .B1(_11523_ ), .B2(_11524_ ), .ZN(_00707_ ) );
NAND4_X1 _15613_ ( .A1(_10371_ ), .A2(_11301_ ), .A3(_11512_ ), .A4(_11493_ ), .ZN(_11525_ ) );
OAI21_X1 _15614_ ( .A(\u_lsu.pmem[3781] ), .B1(_11460_ ), .B2(_10363_ ), .ZN(_11526_ ) );
AOI21_X1 _15615_ ( .A(fanout_net_26 ), .B1(_11525_ ), .B2(_11526_ ), .ZN(_00708_ ) );
OAI21_X1 _15616_ ( .A(\u_lsu.pmem[6534] ), .B1(_11521_ ), .B2(_11522_ ), .ZN(_11527_ ) );
NAND4_X1 _15617_ ( .A1(_09513_ ), .A2(_10185_ ), .A3(_11473_ ), .A4(_11128_ ), .ZN(_11528_ ) );
AOI21_X1 _15618_ ( .A(fanout_net_26 ), .B1(_11527_ ), .B2(_11528_ ), .ZN(_00709_ ) );
OAI21_X1 _15619_ ( .A(\u_lsu.pmem[6533] ), .B1(_11521_ ), .B2(_11522_ ), .ZN(_11529_ ) );
NAND4_X1 _15620_ ( .A1(_09513_ ), .A2(_10188_ ), .A3(_11473_ ), .A4(_11128_ ), .ZN(_11530_ ) );
AOI21_X1 _15621_ ( .A(fanout_net_26 ), .B1(_11529_ ), .B2(_11530_ ), .ZN(_00710_ ) );
OAI21_X1 _15622_ ( .A(\u_lsu.pmem[6532] ), .B1(_11521_ ), .B2(_11522_ ), .ZN(_11531_ ) );
NAND4_X1 _15623_ ( .A1(_09513_ ), .A2(_10192_ ), .A3(_11473_ ), .A4(_11128_ ), .ZN(_11532_ ) );
AOI21_X1 _15624_ ( .A(fanout_net_26 ), .B1(_11531_ ), .B2(_11532_ ), .ZN(_00711_ ) );
OAI21_X1 _15625_ ( .A(\u_lsu.pmem[6531] ), .B1(_11521_ ), .B2(_11522_ ), .ZN(_11533_ ) );
NAND4_X1 _15626_ ( .A1(_09513_ ), .A2(_10915_ ), .A3(_11473_ ), .A4(_11128_ ), .ZN(_11534_ ) );
AOI21_X1 _15627_ ( .A(fanout_net_26 ), .B1(_11533_ ), .B2(_11534_ ), .ZN(_00712_ ) );
OAI21_X1 _15628_ ( .A(\u_lsu.pmem[6530] ), .B1(_11521_ ), .B2(_11522_ ), .ZN(_11535_ ) );
BUF_X4 _15629_ ( .A(_09883_ ), .Z(_11536_ ) );
NAND4_X1 _15630_ ( .A1(_09537_ ), .A2(_11536_ ), .A3(_11473_ ), .A4(_11128_ ), .ZN(_11537_ ) );
AOI21_X1 _15631_ ( .A(fanout_net_26 ), .B1(_11535_ ), .B2(_11537_ ), .ZN(_00713_ ) );
OAI21_X1 _15632_ ( .A(\u_lsu.pmem[6529] ), .B1(_11521_ ), .B2(_11522_ ), .ZN(_11538_ ) );
BUF_X4 _15633_ ( .A(_10904_ ), .Z(_11539_ ) );
NAND4_X1 _15634_ ( .A1(_09513_ ), .A2(_09923_ ), .A3(_11473_ ), .A4(_11539_ ), .ZN(_11540_ ) );
AOI21_X1 _15635_ ( .A(fanout_net_26 ), .B1(_11538_ ), .B2(_11540_ ), .ZN(_00714_ ) );
OAI21_X1 _15636_ ( .A(\u_lsu.pmem[6528] ), .B1(_11521_ ), .B2(_11522_ ), .ZN(_11541_ ) );
BUF_X4 _15637_ ( .A(_09512_ ), .Z(_11542_ ) );
NAND4_X1 _15638_ ( .A1(_11542_ ), .A2(_11131_ ), .A3(_11473_ ), .A4(_11539_ ), .ZN(_11543_ ) );
AOI21_X1 _15639_ ( .A(fanout_net_26 ), .B1(_11541_ ), .B2(_11543_ ), .ZN(_00715_ ) );
NOR2_X1 _15640_ ( .A1(_10397_ ), .A2(_09559_ ), .ZN(_11544_ ) );
AND2_X2 _15641_ ( .A1(_10325_ ), .A2(_11544_ ), .ZN(_11545_ ) );
INV_X1 _15642_ ( .A(_11545_ ), .ZN(_11546_ ) );
BUF_X4 _15643_ ( .A(_11546_ ), .Z(_11547_ ) );
OAI21_X1 _15644_ ( .A(\u_lsu.pmem[6503] ), .B1(_11391_ ), .B2(_11547_ ), .ZN(_11548_ ) );
BUF_X4 _15645_ ( .A(_11545_ ), .Z(_11549_ ) );
NAND3_X1 _15646_ ( .A1(_11138_ ), .A2(_11192_ ), .A3(_11549_ ), .ZN(_11550_ ) );
AOI21_X1 _15647_ ( .A(fanout_net_26 ), .B1(_11548_ ), .B2(_11550_ ), .ZN(_00716_ ) );
OAI21_X1 _15648_ ( .A(\u_lsu.pmem[6502] ), .B1(_11391_ ), .B2(_11547_ ), .ZN(_11551_ ) );
NAND3_X1 _15649_ ( .A1(_10719_ ), .A2(_11192_ ), .A3(_11549_ ), .ZN(_11552_ ) );
AOI21_X1 _15650_ ( .A(fanout_net_26 ), .B1(_11551_ ), .B2(_11552_ ), .ZN(_00717_ ) );
BUF_X4 _15651_ ( .A(_09572_ ), .Z(_11553_ ) );
OAI21_X1 _15652_ ( .A(\u_lsu.pmem[6501] ), .B1(_11553_ ), .B2(_11546_ ), .ZN(_11554_ ) );
NAND3_X1 _15653_ ( .A1(_10728_ ), .A2(_11192_ ), .A3(_11549_ ), .ZN(_11555_ ) );
AOI21_X1 _15654_ ( .A(fanout_net_26 ), .B1(_11554_ ), .B2(_11555_ ), .ZN(_00718_ ) );
NAND4_X1 _15655_ ( .A1(_10374_ ), .A2(_11301_ ), .A3(_11512_ ), .A4(_11493_ ), .ZN(_11556_ ) );
OAI21_X1 _15656_ ( .A(\u_lsu.pmem[3780] ), .B1(_11460_ ), .B2(_10363_ ), .ZN(_11557_ ) );
AOI21_X1 _15657_ ( .A(fanout_net_26 ), .B1(_11556_ ), .B2(_11557_ ), .ZN(_00719_ ) );
OAI21_X1 _15658_ ( .A(\u_lsu.pmem[6500] ), .B1(_11553_ ), .B2(_11546_ ), .ZN(_11558_ ) );
NAND3_X1 _15659_ ( .A1(_11152_ ), .A2(_11192_ ), .A3(_11549_ ), .ZN(_11559_ ) );
AOI21_X1 _15660_ ( .A(fanout_net_26 ), .B1(_11558_ ), .B2(_11559_ ), .ZN(_00720_ ) );
OAI21_X1 _15661_ ( .A(\u_lsu.pmem[6499] ), .B1(_11553_ ), .B2(_11546_ ), .ZN(_11560_ ) );
NAND3_X1 _15662_ ( .A1(_11155_ ), .A2(_11192_ ), .A3(_11549_ ), .ZN(_11561_ ) );
AOI21_X1 _15663_ ( .A(fanout_net_26 ), .B1(_11560_ ), .B2(_11561_ ), .ZN(_00721_ ) );
OAI21_X1 _15664_ ( .A(\u_lsu.pmem[6498] ), .B1(_11553_ ), .B2(_11546_ ), .ZN(_11562_ ) );
NAND3_X1 _15665_ ( .A1(_11158_ ), .A2(_11192_ ), .A3(_11549_ ), .ZN(_11563_ ) );
AOI21_X1 _15666_ ( .A(fanout_net_26 ), .B1(_11562_ ), .B2(_11563_ ), .ZN(_00722_ ) );
OAI21_X1 _15667_ ( .A(\u_lsu.pmem[6497] ), .B1(_11553_ ), .B2(_11546_ ), .ZN(_11564_ ) );
BUF_X4 _15668_ ( .A(_09635_ ), .Z(_11565_ ) );
NAND3_X1 _15669_ ( .A1(_11163_ ), .A2(_11565_ ), .A3(_11549_ ), .ZN(_11566_ ) );
AOI21_X1 _15670_ ( .A(fanout_net_26 ), .B1(_11564_ ), .B2(_11566_ ), .ZN(_00723_ ) );
OAI21_X1 _15671_ ( .A(\u_lsu.pmem[6496] ), .B1(_11553_ ), .B2(_11546_ ), .ZN(_11567_ ) );
NAND3_X1 _15672_ ( .A1(_10741_ ), .A2(_11565_ ), .A3(_11549_ ), .ZN(_11568_ ) );
AOI21_X1 _15673_ ( .A(fanout_net_26 ), .B1(_11567_ ), .B2(_11568_ ), .ZN(_00724_ ) );
NOR2_X1 _15674_ ( .A1(_10397_ ), .A2(_09632_ ), .ZN(_11569_ ) );
AND2_X2 _15675_ ( .A1(_10325_ ), .A2(_11569_ ), .ZN(_11570_ ) );
INV_X1 _15676_ ( .A(_11570_ ), .ZN(_11571_ ) );
BUF_X4 _15677_ ( .A(_11571_ ), .Z(_11572_ ) );
OAI21_X1 _15678_ ( .A(\u_lsu.pmem[6471] ), .B1(_11553_ ), .B2(_11572_ ), .ZN(_11573_ ) );
BUF_X4 _15679_ ( .A(_11570_ ), .Z(_11574_ ) );
NAND3_X1 _15680_ ( .A1(_11138_ ), .A2(_11565_ ), .A3(_11574_ ), .ZN(_11575_ ) );
AOI21_X1 _15681_ ( .A(fanout_net_26 ), .B1(_11573_ ), .B2(_11575_ ), .ZN(_00725_ ) );
OAI21_X1 _15682_ ( .A(\u_lsu.pmem[6470] ), .B1(_11553_ ), .B2(_11572_ ), .ZN(_11576_ ) );
NAND3_X1 _15683_ ( .A1(_10719_ ), .A2(_11565_ ), .A3(_11574_ ), .ZN(_11577_ ) );
AOI21_X1 _15684_ ( .A(fanout_net_26 ), .B1(_11576_ ), .B2(_11577_ ), .ZN(_00726_ ) );
OAI21_X1 _15685_ ( .A(\u_lsu.pmem[6469] ), .B1(_11553_ ), .B2(_11571_ ), .ZN(_11578_ ) );
NAND3_X1 _15686_ ( .A1(_10728_ ), .A2(_11565_ ), .A3(_11574_ ), .ZN(_11579_ ) );
AOI21_X1 _15687_ ( .A(fanout_net_26 ), .B1(_11578_ ), .B2(_11579_ ), .ZN(_00727_ ) );
OAI21_X1 _15688_ ( .A(\u_lsu.pmem[6468] ), .B1(_11553_ ), .B2(_11571_ ), .ZN(_11580_ ) );
NAND3_X1 _15689_ ( .A1(_11152_ ), .A2(_11565_ ), .A3(_11574_ ), .ZN(_11581_ ) );
AOI21_X1 _15690_ ( .A(fanout_net_27 ), .B1(_11580_ ), .B2(_11581_ ), .ZN(_00728_ ) );
BUF_X8 _15691_ ( .A(_09458_ ), .Z(_11582_ ) );
BUF_X4 _15692_ ( .A(_11582_ ), .Z(_11583_ ) );
OAI21_X1 _15693_ ( .A(\u_lsu.pmem[6467] ), .B1(_11583_ ), .B2(_11571_ ), .ZN(_11584_ ) );
NAND3_X1 _15694_ ( .A1(_11155_ ), .A2(_11565_ ), .A3(_11574_ ), .ZN(_11585_ ) );
AOI21_X1 _15695_ ( .A(fanout_net_27 ), .B1(_11584_ ), .B2(_11585_ ), .ZN(_00729_ ) );
NAND4_X1 _15696_ ( .A1(_10377_ ), .A2(_11301_ ), .A3(_11512_ ), .A4(_11493_ ), .ZN(_11586_ ) );
OAI21_X1 _15697_ ( .A(\u_lsu.pmem[3779] ), .B1(_11460_ ), .B2(_10363_ ), .ZN(_11587_ ) );
AOI21_X1 _15698_ ( .A(fanout_net_27 ), .B1(_11586_ ), .B2(_11587_ ), .ZN(_00730_ ) );
OAI21_X1 _15699_ ( .A(\u_lsu.pmem[6466] ), .B1(_11583_ ), .B2(_11571_ ), .ZN(_11588_ ) );
NAND3_X1 _15700_ ( .A1(_11158_ ), .A2(_11565_ ), .A3(_11574_ ), .ZN(_11589_ ) );
AOI21_X1 _15701_ ( .A(fanout_net_27 ), .B1(_11588_ ), .B2(_11589_ ), .ZN(_00731_ ) );
OAI21_X1 _15702_ ( .A(\u_lsu.pmem[6465] ), .B1(_11583_ ), .B2(_11571_ ), .ZN(_11590_ ) );
NAND3_X1 _15703_ ( .A1(_11163_ ), .A2(_11565_ ), .A3(_11574_ ), .ZN(_11591_ ) );
AOI21_X1 _15704_ ( .A(fanout_net_27 ), .B1(_11590_ ), .B2(_11591_ ), .ZN(_00732_ ) );
OAI21_X1 _15705_ ( .A(\u_lsu.pmem[6464] ), .B1(_11583_ ), .B2(_11571_ ), .ZN(_11592_ ) );
NAND3_X1 _15706_ ( .A1(_10741_ ), .A2(_11565_ ), .A3(_11574_ ), .ZN(_11593_ ) );
AOI21_X1 _15707_ ( .A(fanout_net_27 ), .B1(_11592_ ), .B2(_11593_ ), .ZN(_00733_ ) );
BUF_X4 _15708_ ( .A(_11453_ ), .Z(_11594_ ) );
NAND4_X1 _15709_ ( .A1(_09670_ ), .A2(_11594_ ), .A3(_11512_ ), .A4(_11515_ ), .ZN(_11595_ ) );
AND2_X2 _15710_ ( .A1(_09131_ ), .A2(_09135_ ), .ZN(_11596_ ) );
INV_X1 _15711_ ( .A(_11596_ ), .ZN(_11597_ ) );
BUF_X4 _15712_ ( .A(_11597_ ), .Z(_11598_ ) );
OAI21_X1 _15713_ ( .A(\u_lsu.pmem[6439] ), .B1(_11598_ ), .B2(_11337_ ), .ZN(_11599_ ) );
AOI21_X1 _15714_ ( .A(fanout_net_27 ), .B1(_11595_ ), .B2(_11599_ ), .ZN(_00734_ ) );
NAND4_X1 _15715_ ( .A1(_09681_ ), .A2(_11594_ ), .A3(_11512_ ), .A4(_11515_ ), .ZN(_11600_ ) );
OAI21_X1 _15716_ ( .A(\u_lsu.pmem[6438] ), .B1(_11598_ ), .B2(_11337_ ), .ZN(_11601_ ) );
AOI21_X1 _15717_ ( .A(fanout_net_27 ), .B1(_11600_ ), .B2(_11601_ ), .ZN(_00735_ ) );
NAND4_X1 _15718_ ( .A1(_09685_ ), .A2(_11594_ ), .A3(_11512_ ), .A4(_11515_ ), .ZN(_11602_ ) );
OAI21_X1 _15719_ ( .A(\u_lsu.pmem[6437] ), .B1(_11598_ ), .B2(_11337_ ), .ZN(_11603_ ) );
AOI21_X1 _15720_ ( .A(fanout_net_27 ), .B1(_11602_ ), .B2(_11603_ ), .ZN(_00736_ ) );
AND2_X1 _15721_ ( .A1(_11596_ ), .A2(_09141_ ), .ZN(_11604_ ) );
OAI21_X1 _15722_ ( .A(_10715_ ), .B1(_11604_ ), .B2(\u_lsu.pmem[6436] ), .ZN(_11605_ ) );
AOI21_X1 _15723_ ( .A(_11605_ ), .B1(_09691_ ), .B2(_11604_ ), .ZN(_00737_ ) );
OAI21_X1 _15724_ ( .A(\u_lsu.pmem[6435] ), .B1(_11598_ ), .B2(_11522_ ), .ZN(_11606_ ) );
NAND3_X1 _15725_ ( .A1(_10733_ ), .A2(_11596_ ), .A3(_11426_ ), .ZN(_11607_ ) );
AOI21_X1 _15726_ ( .A(fanout_net_27 ), .B1(_11606_ ), .B2(_11607_ ), .ZN(_00738_ ) );
OAI21_X1 _15727_ ( .A(\u_lsu.pmem[6434] ), .B1(_11598_ ), .B2(_11522_ ), .ZN(_02187_ ) );
NAND3_X1 _15728_ ( .A1(_11158_ ), .A2(_11596_ ), .A3(_11426_ ), .ZN(_02188_ ) );
AOI21_X1 _15729_ ( .A(fanout_net_27 ), .B1(_02187_ ), .B2(_02188_ ), .ZN(_00739_ ) );
BUF_X4 _15730_ ( .A(_10901_ ), .Z(_02189_ ) );
OAI21_X1 _15731_ ( .A(\u_lsu.pmem[6433] ), .B1(_11598_ ), .B2(_02189_ ), .ZN(_02190_ ) );
NAND3_X1 _15732_ ( .A1(_10738_ ), .A2(_11596_ ), .A3(_11426_ ), .ZN(_02191_ ) );
AOI21_X1 _15733_ ( .A(fanout_net_27 ), .B1(_02190_ ), .B2(_02191_ ), .ZN(_00740_ ) );
NAND4_X1 _15734_ ( .A1(_10381_ ), .A2(_11301_ ), .A3(_11512_ ), .A4(_11493_ ), .ZN(_02192_ ) );
OAI21_X1 _15735_ ( .A(\u_lsu.pmem[3778] ), .B1(_11460_ ), .B2(_10363_ ), .ZN(_02193_ ) );
AOI21_X1 _15736_ ( .A(fanout_net_27 ), .B1(_02192_ ), .B2(_02193_ ), .ZN(_00741_ ) );
NAND4_X1 _15737_ ( .A1(_09703_ ), .A2(_11594_ ), .A3(_11512_ ), .A4(_11515_ ), .ZN(_02194_ ) );
OAI21_X1 _15738_ ( .A(\u_lsu.pmem[6432] ), .B1(_11598_ ), .B2(_11337_ ), .ZN(_02195_ ) );
AOI21_X1 _15739_ ( .A(fanout_net_27 ), .B1(_02194_ ), .B2(_02195_ ), .ZN(_00742_ ) );
BUF_X8 _15740_ ( .A(_09877_ ), .Z(_02196_ ) );
BUF_X4 _15741_ ( .A(_02196_ ), .Z(_02197_ ) );
NAND4_X1 _15742_ ( .A1(_09708_ ), .A2(_11594_ ), .A3(_02197_ ), .A4(_11515_ ), .ZN(_02198_ ) );
NAND2_X1 _15743_ ( .A1(_09467_ ), .A2(_10424_ ), .ZN(_02199_ ) );
BUF_X4 _15744_ ( .A(_02199_ ), .Z(_02200_ ) );
OAI21_X1 _15745_ ( .A(\u_lsu.pmem[6407] ), .B1(_11504_ ), .B2(_02200_ ), .ZN(_02201_ ) );
AOI21_X1 _15746_ ( .A(fanout_net_27 ), .B1(_02198_ ), .B2(_02201_ ), .ZN(_00743_ ) );
NAND4_X1 _15747_ ( .A1(_09715_ ), .A2(_11594_ ), .A3(_02197_ ), .A4(_11515_ ), .ZN(_02202_ ) );
OAI21_X1 _15748_ ( .A(\u_lsu.pmem[6406] ), .B1(_11504_ ), .B2(_02200_ ), .ZN(_02203_ ) );
AOI21_X1 _15749_ ( .A(fanout_net_27 ), .B1(_02202_ ), .B2(_02203_ ), .ZN(_00744_ ) );
NAND4_X1 _15750_ ( .A1(_09718_ ), .A2(_11594_ ), .A3(_02197_ ), .A4(_11515_ ), .ZN(_02204_ ) );
OAI21_X1 _15751_ ( .A(\u_lsu.pmem[6405] ), .B1(_11504_ ), .B2(_02200_ ), .ZN(_02205_ ) );
AOI21_X1 _15752_ ( .A(fanout_net_27 ), .B1(_02204_ ), .B2(_02205_ ), .ZN(_00745_ ) );
NAND4_X1 _15753_ ( .A1(_09721_ ), .A2(_11594_ ), .A3(_02197_ ), .A4(_11515_ ), .ZN(_02206_ ) );
OAI21_X1 _15754_ ( .A(\u_lsu.pmem[6404] ), .B1(_11504_ ), .B2(_02200_ ), .ZN(_02207_ ) );
AOI21_X1 _15755_ ( .A(fanout_net_27 ), .B1(_02206_ ), .B2(_02207_ ), .ZN(_00746_ ) );
NAND4_X1 _15756_ ( .A1(_09725_ ), .A2(_11594_ ), .A3(_02197_ ), .A4(_11515_ ), .ZN(_02208_ ) );
BUF_X8 _15757_ ( .A(_09458_ ), .Z(_02209_ ) );
BUF_X4 _15758_ ( .A(_02209_ ), .Z(_02210_ ) );
OAI21_X1 _15759_ ( .A(\u_lsu.pmem[6403] ), .B1(_02210_ ), .B2(_02200_ ), .ZN(_02211_ ) );
AOI21_X1 _15760_ ( .A(fanout_net_27 ), .B1(_02208_ ), .B2(_02211_ ), .ZN(_00747_ ) );
OAI21_X1 _15761_ ( .A(\u_lsu.pmem[6402] ), .B1(_11583_ ), .B2(_02200_ ), .ZN(_02212_ ) );
BUF_X4 _15762_ ( .A(_11381_ ), .Z(_02213_ ) );
NAND4_X1 _15763_ ( .A1(_09510_ ), .A2(_09474_ ), .A3(_02213_ ), .A4(_09467_ ), .ZN(_02214_ ) );
AOI21_X1 _15764_ ( .A(fanout_net_27 ), .B1(_02212_ ), .B2(_02214_ ), .ZN(_00748_ ) );
BUF_X4 _15765_ ( .A(_11334_ ), .Z(_02215_ ) );
NAND4_X1 _15766_ ( .A1(_09733_ ), .A2(_11594_ ), .A3(_02197_ ), .A4(_02215_ ), .ZN(_02216_ ) );
OAI21_X1 _15767_ ( .A(\u_lsu.pmem[6401] ), .B1(_02210_ ), .B2(_02200_ ), .ZN(_02217_ ) );
AOI21_X1 _15768_ ( .A(fanout_net_27 ), .B1(_02216_ ), .B2(_02217_ ), .ZN(_00749_ ) );
BUF_X4 _15769_ ( .A(_11453_ ), .Z(_02218_ ) );
NAND4_X1 _15770_ ( .A1(_09736_ ), .A2(_02218_ ), .A3(_02197_ ), .A4(_02215_ ), .ZN(_02219_ ) );
OAI21_X1 _15771_ ( .A(\u_lsu.pmem[6400] ), .B1(_02210_ ), .B2(_02200_ ), .ZN(_02220_ ) );
AOI21_X1 _15772_ ( .A(fanout_net_27 ), .B1(_02219_ ), .B2(_02220_ ), .ZN(_00750_ ) );
NAND2_X4 _15773_ ( .A1(_11028_ ), .A2(_09749_ ), .ZN(_02221_ ) );
BUF_X4 _15774_ ( .A(_02221_ ), .Z(_02222_ ) );
OAI21_X1 _15775_ ( .A(\u_lsu.pmem[6375] ), .B1(_11583_ ), .B2(_02222_ ), .ZN(_02223_ ) );
NAND4_X1 _15776_ ( .A1(_10851_ ), .A2(_11393_ ), .A3(_02213_ ), .A4(_09749_ ), .ZN(_02224_ ) );
AOI21_X1 _15777_ ( .A(fanout_net_27 ), .B1(_02223_ ), .B2(_02224_ ), .ZN(_00751_ ) );
BUF_X4 _15778_ ( .A(_10886_ ), .Z(_02225_ ) );
NAND4_X1 _15779_ ( .A1(_10384_ ), .A2(_02225_ ), .A3(_02197_ ), .A4(_11493_ ), .ZN(_02226_ ) );
OAI21_X1 _15780_ ( .A(\u_lsu.pmem[3777] ), .B1(_11460_ ), .B2(_10363_ ), .ZN(_02227_ ) );
AOI21_X1 _15781_ ( .A(fanout_net_27 ), .B1(_02226_ ), .B2(_02227_ ), .ZN(_00752_ ) );
NAND4_X1 _15782_ ( .A1(_09756_ ), .A2(_02218_ ), .A3(_02197_ ), .A4(_02215_ ), .ZN(_02228_ ) );
OAI21_X1 _15783_ ( .A(\u_lsu.pmem[6374] ), .B1(_02210_ ), .B2(_02222_ ), .ZN(_02229_ ) );
AOI21_X1 _15784_ ( .A(fanout_net_27 ), .B1(_02228_ ), .B2(_02229_ ), .ZN(_00753_ ) );
NAND4_X1 _15785_ ( .A1(_09763_ ), .A2(_02218_ ), .A3(_02197_ ), .A4(_02215_ ), .ZN(_02230_ ) );
OAI21_X1 _15786_ ( .A(\u_lsu.pmem[6373] ), .B1(_02210_ ), .B2(_02222_ ), .ZN(_02231_ ) );
AOI21_X1 _15787_ ( .A(fanout_net_27 ), .B1(_02230_ ), .B2(_02231_ ), .ZN(_00754_ ) );
BUF_X4 _15788_ ( .A(_02196_ ), .Z(_02232_ ) );
NAND4_X1 _15789_ ( .A1(_09770_ ), .A2(_02218_ ), .A3(_02232_ ), .A4(_02215_ ), .ZN(_02233_ ) );
OAI21_X1 _15790_ ( .A(\u_lsu.pmem[6372] ), .B1(_02210_ ), .B2(_02222_ ), .ZN(_02234_ ) );
AOI21_X1 _15791_ ( .A(fanout_net_27 ), .B1(_02233_ ), .B2(_02234_ ), .ZN(_00755_ ) );
NAND4_X1 _15792_ ( .A1(_09775_ ), .A2(_02218_ ), .A3(_02232_ ), .A4(_02215_ ), .ZN(_02235_ ) );
OAI21_X1 _15793_ ( .A(\u_lsu.pmem[6371] ), .B1(_02210_ ), .B2(_02222_ ), .ZN(_02236_ ) );
AOI21_X1 _15794_ ( .A(fanout_net_27 ), .B1(_02235_ ), .B2(_02236_ ), .ZN(_00756_ ) );
NAND4_X1 _15795_ ( .A1(_09780_ ), .A2(_02218_ ), .A3(_02232_ ), .A4(_02215_ ), .ZN(_02237_ ) );
OAI21_X1 _15796_ ( .A(\u_lsu.pmem[6370] ), .B1(_02210_ ), .B2(_02222_ ), .ZN(_02238_ ) );
AOI21_X1 _15797_ ( .A(fanout_net_27 ), .B1(_02237_ ), .B2(_02238_ ), .ZN(_00757_ ) );
NAND4_X1 _15798_ ( .A1(_09787_ ), .A2(_02218_ ), .A3(_02232_ ), .A4(_02215_ ), .ZN(_02239_ ) );
OAI21_X1 _15799_ ( .A(\u_lsu.pmem[6369] ), .B1(_02210_ ), .B2(_02222_ ), .ZN(_02240_ ) );
AOI21_X1 _15800_ ( .A(fanout_net_27 ), .B1(_02239_ ), .B2(_02240_ ), .ZN(_00758_ ) );
NAND4_X1 _15801_ ( .A1(_09791_ ), .A2(_02218_ ), .A3(_02232_ ), .A4(_02215_ ), .ZN(_02241_ ) );
OAI21_X1 _15802_ ( .A(\u_lsu.pmem[6368] ), .B1(_02210_ ), .B2(_02222_ ), .ZN(_02242_ ) );
AOI21_X1 _15803_ ( .A(fanout_net_28 ), .B1(_02241_ ), .B2(_02242_ ), .ZN(_00759_ ) );
NAND2_X4 _15804_ ( .A1(_11028_ ), .A2(_09798_ ), .ZN(_02243_ ) );
BUF_X4 _15805_ ( .A(_02243_ ), .Z(_02244_ ) );
OAI21_X1 _15806_ ( .A(\u_lsu.pmem[6343] ), .B1(_11583_ ), .B2(_02244_ ), .ZN(_02245_ ) );
BUF_X4 _15807_ ( .A(_09741_ ), .Z(_02246_ ) );
NAND4_X1 _15808_ ( .A1(_02246_ ), .A2(_11393_ ), .A3(_02213_ ), .A4(_09798_ ), .ZN(_02247_ ) );
AOI21_X1 _15809_ ( .A(fanout_net_28 ), .B1(_02245_ ), .B2(_02247_ ), .ZN(_00760_ ) );
NAND4_X1 _15810_ ( .A1(_09804_ ), .A2(_09806_ ), .A3(_02232_ ), .A4(_02215_ ), .ZN(_02248_ ) );
BUF_X4 _15811_ ( .A(_02209_ ), .Z(_02249_ ) );
OAI21_X1 _15812_ ( .A(\u_lsu.pmem[6342] ), .B1(_02249_ ), .B2(_02244_ ), .ZN(_02250_ ) );
AOI21_X1 _15813_ ( .A(fanout_net_28 ), .B1(_02248_ ), .B2(_02250_ ), .ZN(_00761_ ) );
BUF_X4 _15814_ ( .A(_11334_ ), .Z(_02251_ ) );
NAND4_X1 _15815_ ( .A1(_09811_ ), .A2(_02218_ ), .A3(_02232_ ), .A4(_02251_ ), .ZN(_02252_ ) );
OAI21_X1 _15816_ ( .A(\u_lsu.pmem[6341] ), .B1(_02249_ ), .B2(_02244_ ), .ZN(_02253_ ) );
AOI21_X1 _15817_ ( .A(fanout_net_28 ), .B1(_02252_ ), .B2(_02253_ ), .ZN(_00762_ ) );
NAND4_X1 _15818_ ( .A1(_10391_ ), .A2(_02225_ ), .A3(_02232_ ), .A4(_11493_ ), .ZN(_02254_ ) );
OAI21_X1 _15819_ ( .A(\u_lsu.pmem[3776] ), .B1(_11460_ ), .B2(_10363_ ), .ZN(_02255_ ) );
AOI21_X1 _15820_ ( .A(fanout_net_28 ), .B1(_02254_ ), .B2(_02255_ ), .ZN(_00763_ ) );
NAND4_X1 _15821_ ( .A1(_09815_ ), .A2(_02218_ ), .A3(_02232_ ), .A4(_02251_ ), .ZN(_02256_ ) );
OAI21_X1 _15822_ ( .A(\u_lsu.pmem[6340] ), .B1(_02249_ ), .B2(_02244_ ), .ZN(_02257_ ) );
AOI21_X1 _15823_ ( .A(fanout_net_28 ), .B1(_02256_ ), .B2(_02257_ ), .ZN(_00764_ ) );
BUF_X4 _15824_ ( .A(_11453_ ), .Z(_02258_ ) );
NAND4_X1 _15825_ ( .A1(_09819_ ), .A2(_02258_ ), .A3(_02232_ ), .A4(_02251_ ), .ZN(_02259_ ) );
OAI21_X1 _15826_ ( .A(\u_lsu.pmem[6339] ), .B1(_02249_ ), .B2(_02244_ ), .ZN(_02260_ ) );
AOI21_X1 _15827_ ( .A(fanout_net_28 ), .B1(_02259_ ), .B2(_02260_ ), .ZN(_00765_ ) );
BUF_X4 _15828_ ( .A(_02196_ ), .Z(_02261_ ) );
NAND4_X1 _15829_ ( .A1(_09827_ ), .A2(_02258_ ), .A3(_02261_ ), .A4(_02251_ ), .ZN(_02262_ ) );
OAI21_X1 _15830_ ( .A(\u_lsu.pmem[6338] ), .B1(_02249_ ), .B2(_02244_ ), .ZN(_02263_ ) );
AOI21_X1 _15831_ ( .A(fanout_net_28 ), .B1(_02262_ ), .B2(_02263_ ), .ZN(_00766_ ) );
NAND4_X1 _15832_ ( .A1(_09831_ ), .A2(_02258_ ), .A3(_02261_ ), .A4(_02251_ ), .ZN(_02264_ ) );
OAI21_X1 _15833_ ( .A(\u_lsu.pmem[6337] ), .B1(_02249_ ), .B2(_02244_ ), .ZN(_02265_ ) );
AOI21_X1 _15834_ ( .A(fanout_net_28 ), .B1(_02264_ ), .B2(_02265_ ), .ZN(_00767_ ) );
NAND4_X1 _15835_ ( .A1(_09835_ ), .A2(_02258_ ), .A3(_02261_ ), .A4(_02251_ ), .ZN(_02266_ ) );
OAI21_X1 _15836_ ( .A(\u_lsu.pmem[6336] ), .B1(_02249_ ), .B2(_02244_ ), .ZN(_02267_ ) );
AOI21_X1 _15837_ ( .A(fanout_net_28 ), .B1(_02266_ ), .B2(_02267_ ), .ZN(_00768_ ) );
NAND4_X1 _15838_ ( .A1(_09840_ ), .A2(_02258_ ), .A3(_02261_ ), .A4(_02251_ ), .ZN(_02268_ ) );
NAND3_X1 _15839_ ( .A1(_10424_ ), .A2(_09842_ ), .A3(_09844_ ), .ZN(_02269_ ) );
BUF_X4 _15840_ ( .A(_02269_ ), .Z(_02270_ ) );
OAI21_X1 _15841_ ( .A(\u_lsu.pmem[6311] ), .B1(_02249_ ), .B2(_02270_ ), .ZN(_02271_ ) );
AOI21_X1 _15842_ ( .A(fanout_net_28 ), .B1(_02268_ ), .B2(_02271_ ), .ZN(_00769_ ) );
NAND4_X1 _15843_ ( .A1(_09849_ ), .A2(_02258_ ), .A3(_02261_ ), .A4(_02251_ ), .ZN(_02272_ ) );
OAI21_X1 _15844_ ( .A(\u_lsu.pmem[6310] ), .B1(_02249_ ), .B2(_02270_ ), .ZN(_02273_ ) );
AOI21_X1 _15845_ ( .A(fanout_net_28 ), .B1(_02272_ ), .B2(_02273_ ), .ZN(_00770_ ) );
NAND4_X1 _15846_ ( .A1(_09853_ ), .A2(_02258_ ), .A3(_02261_ ), .A4(_02251_ ), .ZN(_02274_ ) );
OAI21_X1 _15847_ ( .A(\u_lsu.pmem[6309] ), .B1(_02249_ ), .B2(_02270_ ), .ZN(_02275_ ) );
AOI21_X1 _15848_ ( .A(fanout_net_28 ), .B1(_02274_ ), .B2(_02275_ ), .ZN(_00771_ ) );
NAND4_X1 _15849_ ( .A1(_09858_ ), .A2(_02258_ ), .A3(_02261_ ), .A4(_02251_ ), .ZN(_02276_ ) );
BUF_X4 _15850_ ( .A(_02209_ ), .Z(_02277_ ) );
OAI21_X1 _15851_ ( .A(\u_lsu.pmem[6308] ), .B1(_02277_ ), .B2(_02270_ ), .ZN(_02278_ ) );
AOI21_X1 _15852_ ( .A(fanout_net_28 ), .B1(_02276_ ), .B2(_02278_ ), .ZN(_00772_ ) );
BUF_X4 _15853_ ( .A(_11334_ ), .Z(_02279_ ) );
NAND4_X1 _15854_ ( .A1(_09861_ ), .A2(_02258_ ), .A3(_02261_ ), .A4(_02279_ ), .ZN(_02280_ ) );
OAI21_X1 _15855_ ( .A(\u_lsu.pmem[6307] ), .B1(_02277_ ), .B2(_02270_ ), .ZN(_02281_ ) );
AOI21_X1 _15856_ ( .A(fanout_net_28 ), .B1(_02280_ ), .B2(_02281_ ), .ZN(_00773_ ) );
NAND4_X1 _15857_ ( .A1(_10394_ ), .A2(_02225_ ), .A3(_02261_ ), .A4(_11493_ ), .ZN(_02282_ ) );
OAI21_X1 _15858_ ( .A(\u_lsu.pmem[3751] ), .B1(_11460_ ), .B2(_10400_ ), .ZN(_02283_ ) );
AOI21_X1 _15859_ ( .A(fanout_net_28 ), .B1(_02282_ ), .B2(_02283_ ), .ZN(_00774_ ) );
NAND4_X1 _15860_ ( .A1(_09864_ ), .A2(_02258_ ), .A3(_02261_ ), .A4(_02279_ ), .ZN(_02284_ ) );
OAI21_X1 _15861_ ( .A(\u_lsu.pmem[6306] ), .B1(_02277_ ), .B2(_02270_ ), .ZN(_02285_ ) );
AOI21_X1 _15862_ ( .A(fanout_net_28 ), .B1(_02284_ ), .B2(_02285_ ), .ZN(_00775_ ) );
BUF_X4 _15863_ ( .A(_11453_ ), .Z(_02286_ ) );
BUF_X4 _15864_ ( .A(_02196_ ), .Z(_02287_ ) );
NAND4_X1 _15865_ ( .A1(_09867_ ), .A2(_02286_ ), .A3(_02287_ ), .A4(_02279_ ), .ZN(_02288_ ) );
OAI21_X1 _15866_ ( .A(\u_lsu.pmem[6305] ), .B1(_02277_ ), .B2(_02270_ ), .ZN(_02289_ ) );
AOI21_X1 _15867_ ( .A(fanout_net_28 ), .B1(_02288_ ), .B2(_02289_ ), .ZN(_00776_ ) );
NAND4_X1 _15868_ ( .A1(_09881_ ), .A2(_02286_ ), .A3(_02287_ ), .A4(_02279_ ), .ZN(_02290_ ) );
OAI21_X1 _15869_ ( .A(\u_lsu.pmem[6304] ), .B1(_02277_ ), .B2(_02270_ ), .ZN(_02291_ ) );
AOI21_X1 _15870_ ( .A(fanout_net_28 ), .B1(_02290_ ), .B2(_02291_ ), .ZN(_00777_ ) );
OR3_X4 _15871_ ( .A1(_09889_ ), .A2(_09743_ ), .A3(_09454_ ), .ZN(_02292_ ) );
BUF_X4 _15872_ ( .A(_02292_ ), .Z(_02293_ ) );
OAI21_X1 _15873_ ( .A(\u_lsu.pmem[6279] ), .B1(_02293_ ), .B2(_02189_ ), .ZN(_02294_ ) );
NAND4_X1 _15874_ ( .A1(_09894_ ), .A2(_10752_ ), .A3(_02213_ ), .A4(_11539_ ), .ZN(_02295_ ) );
AOI21_X1 _15875_ ( .A(fanout_net_28 ), .B1(_02294_ ), .B2(_02295_ ), .ZN(_00778_ ) );
OAI21_X1 _15876_ ( .A(\u_lsu.pmem[6278] ), .B1(_02293_ ), .B2(_02189_ ), .ZN(_02296_ ) );
NAND4_X1 _15877_ ( .A1(_09894_ ), .A2(_10185_ ), .A3(_02213_ ), .A4(_11539_ ), .ZN(_02297_ ) );
AOI21_X1 _15878_ ( .A(fanout_net_28 ), .B1(_02296_ ), .B2(_02297_ ), .ZN(_00779_ ) );
OAI21_X1 _15879_ ( .A(\u_lsu.pmem[6277] ), .B1(_02293_ ), .B2(_02189_ ), .ZN(_02298_ ) );
NAND4_X1 _15880_ ( .A1(_09894_ ), .A2(_10188_ ), .A3(_02213_ ), .A4(_11539_ ), .ZN(_02299_ ) );
AOI21_X1 _15881_ ( .A(fanout_net_28 ), .B1(_02298_ ), .B2(_02299_ ), .ZN(_00780_ ) );
OAI21_X1 _15882_ ( .A(\u_lsu.pmem[6276] ), .B1(_02293_ ), .B2(_02189_ ), .ZN(_02300_ ) );
BUF_X4 _15883_ ( .A(_09893_ ), .Z(_02301_ ) );
NAND4_X1 _15884_ ( .A1(_02301_ ), .A2(_10192_ ), .A3(_02213_ ), .A4(_11539_ ), .ZN(_02302_ ) );
AOI21_X1 _15885_ ( .A(fanout_net_28 ), .B1(_02300_ ), .B2(_02302_ ), .ZN(_00781_ ) );
OAI21_X1 _15886_ ( .A(\u_lsu.pmem[6275] ), .B1(_02293_ ), .B2(_02189_ ), .ZN(_02303_ ) );
NAND4_X1 _15887_ ( .A1(_02301_ ), .A2(_10915_ ), .A3(_02213_ ), .A4(_11539_ ), .ZN(_02304_ ) );
AOI21_X1 _15888_ ( .A(fanout_net_28 ), .B1(_02303_ ), .B2(_02304_ ), .ZN(_00782_ ) );
OAI21_X1 _15889_ ( .A(\u_lsu.pmem[6274] ), .B1(_02293_ ), .B2(_02189_ ), .ZN(_02305_ ) );
NAND4_X1 _15890_ ( .A1(_09906_ ), .A2(_11536_ ), .A3(_02213_ ), .A4(_11539_ ), .ZN(_02306_ ) );
AOI21_X1 _15891_ ( .A(fanout_net_28 ), .B1(_02305_ ), .B2(_02306_ ), .ZN(_00783_ ) );
OAI21_X1 _15892_ ( .A(\u_lsu.pmem[6273] ), .B1(_02293_ ), .B2(_02189_ ), .ZN(_02307_ ) );
BUF_X4 _15893_ ( .A(_09543_ ), .Z(_02308_ ) );
NAND4_X1 _15894_ ( .A1(_02301_ ), .A2(_02308_ ), .A3(_02213_ ), .A4(_11539_ ), .ZN(_02309_ ) );
AOI21_X1 _15895_ ( .A(fanout_net_28 ), .B1(_02307_ ), .B2(_02309_ ), .ZN(_00784_ ) );
NAND4_X1 _15896_ ( .A1(_10402_ ), .A2(_02225_ ), .A3(_02287_ ), .A4(_11493_ ), .ZN(_02310_ ) );
OAI21_X1 _15897_ ( .A(\u_lsu.pmem[3750] ), .B1(_11460_ ), .B2(_10400_ ), .ZN(_02311_ ) );
AOI21_X1 _15898_ ( .A(fanout_net_28 ), .B1(_02310_ ), .B2(_02311_ ), .ZN(_00785_ ) );
OAI21_X1 _15899_ ( .A(\u_lsu.pmem[6272] ), .B1(_02293_ ), .B2(_02189_ ), .ZN(_02312_ ) );
BUF_X4 _15900_ ( .A(_11381_ ), .Z(_02313_ ) );
NAND4_X1 _15901_ ( .A1(_02301_ ), .A2(_11131_ ), .A3(_02313_ ), .A4(_11539_ ), .ZN(_02314_ ) );
AOI21_X1 _15902_ ( .A(fanout_net_28 ), .B1(_02312_ ), .B2(_02314_ ), .ZN(_00786_ ) );
NAND3_X1 _15903_ ( .A1(_09134_ ), .A2(_09506_ ), .A3(_09915_ ), .ZN(_02315_ ) );
BUF_X4 _15904_ ( .A(_02315_ ), .Z(_02316_ ) );
OAI21_X1 _15905_ ( .A(\u_lsu.pmem[6247] ), .B1(_11583_ ), .B2(_02316_ ), .ZN(_02317_ ) );
BUF_X4 _15906_ ( .A(_10548_ ), .Z(_02318_ ) );
NAND4_X1 _15907_ ( .A1(_02246_ ), .A2(_02318_ ), .A3(_02313_ ), .A4(_09917_ ), .ZN(_02319_ ) );
AOI21_X1 _15908_ ( .A(fanout_net_28 ), .B1(_02317_ ), .B2(_02319_ ), .ZN(_00787_ ) );
OAI21_X1 _15909_ ( .A(\u_lsu.pmem[6246] ), .B1(_11583_ ), .B2(_02316_ ), .ZN(_02320_ ) );
NAND4_X1 _15910_ ( .A1(_11347_ ), .A2(_02318_ ), .A3(_02313_ ), .A4(_09917_ ), .ZN(_02321_ ) );
AOI21_X1 _15911_ ( .A(fanout_net_28 ), .B1(_02320_ ), .B2(_02321_ ), .ZN(_00788_ ) );
OAI21_X1 _15912_ ( .A(\u_lsu.pmem[6245] ), .B1(_11583_ ), .B2(_02316_ ), .ZN(_02322_ ) );
BUF_X4 _15913_ ( .A(_09916_ ), .Z(_02323_ ) );
NAND4_X1 _15914_ ( .A1(_11351_ ), .A2(_02318_ ), .A3(_02313_ ), .A4(_02323_ ), .ZN(_02324_ ) );
AOI21_X1 _15915_ ( .A(fanout_net_29 ), .B1(_02322_ ), .B2(_02324_ ), .ZN(_00789_ ) );
BUF_X4 _15916_ ( .A(_11582_ ), .Z(_02325_ ) );
OAI21_X1 _15917_ ( .A(\u_lsu.pmem[6244] ), .B1(_02325_ ), .B2(_02316_ ), .ZN(_02326_ ) );
BUF_X4 _15918_ ( .A(_09148_ ), .Z(_02327_ ) );
NAND4_X1 _15919_ ( .A1(_02327_ ), .A2(_02318_ ), .A3(_02313_ ), .A4(_02323_ ), .ZN(_02328_ ) );
AOI21_X1 _15920_ ( .A(fanout_net_29 ), .B1(_02326_ ), .B2(_02328_ ), .ZN(_00790_ ) );
OAI21_X1 _15921_ ( .A(\u_lsu.pmem[6243] ), .B1(_02325_ ), .B2(_02316_ ), .ZN(_02329_ ) );
NAND4_X1 _15922_ ( .A1(_11385_ ), .A2(_02318_ ), .A3(_02313_ ), .A4(_02323_ ), .ZN(_02330_ ) );
AOI21_X1 _15923_ ( .A(fanout_net_29 ), .B1(_02329_ ), .B2(_02330_ ), .ZN(_00791_ ) );
OAI21_X1 _15924_ ( .A(\u_lsu.pmem[6242] ), .B1(_02325_ ), .B2(_02316_ ), .ZN(_02331_ ) );
NAND4_X1 _15925_ ( .A1(_10492_ ), .A2(_02318_ ), .A3(_02313_ ), .A4(_02323_ ), .ZN(_02332_ ) );
AOI21_X1 _15926_ ( .A(fanout_net_29 ), .B1(_02331_ ), .B2(_02332_ ), .ZN(_00792_ ) );
OAI21_X1 _15927_ ( .A(\u_lsu.pmem[6241] ), .B1(_02325_ ), .B2(_02316_ ), .ZN(_02333_ ) );
NAND4_X1 _15928_ ( .A1(_11414_ ), .A2(_02318_ ), .A3(_02313_ ), .A4(_02323_ ), .ZN(_02334_ ) );
AOI21_X1 _15929_ ( .A(fanout_net_29 ), .B1(_02333_ ), .B2(_02334_ ), .ZN(_00793_ ) );
OAI21_X1 _15930_ ( .A(\u_lsu.pmem[6240] ), .B1(_02325_ ), .B2(_02316_ ), .ZN(_02335_ ) );
NAND4_X1 _15931_ ( .A1(_10525_ ), .A2(_02318_ ), .A3(_02313_ ), .A4(_02323_ ), .ZN(_02336_ ) );
AOI21_X1 _15932_ ( .A(fanout_net_29 ), .B1(_02335_ ), .B2(_02336_ ), .ZN(_00794_ ) );
NAND3_X4 _15933_ ( .A1(_09135_ ), .A2(_09842_ ), .A3(_09948_ ), .ZN(_02337_ ) );
OR4_X2 _15934_ ( .A1(_09565_ ), .A2(_02337_ ), .A3(_11011_ ), .A4(_10873_ ), .ZN(_02338_ ) );
BUF_X4 _15935_ ( .A(_02337_ ), .Z(_02339_ ) );
OAI21_X1 _15936_ ( .A(\u_lsu.pmem[6215] ), .B1(_02277_ ), .B2(_02339_ ), .ZN(_02340_ ) );
AOI21_X1 _15937_ ( .A(fanout_net_29 ), .B1(_02338_ ), .B2(_02340_ ), .ZN(_00795_ ) );
NAND4_X1 _15938_ ( .A1(_10405_ ), .A2(_02225_ ), .A3(_02287_ ), .A4(_11493_ ), .ZN(_02341_ ) );
BUF_X4 _15939_ ( .A(_09562_ ), .Z(_02342_ ) );
OAI21_X1 _15940_ ( .A(\u_lsu.pmem[3749] ), .B1(_02342_ ), .B2(_10399_ ), .ZN(_02343_ ) );
AOI21_X1 _15941_ ( .A(fanout_net_29 ), .B1(_02341_ ), .B2(_02343_ ), .ZN(_00796_ ) );
OAI21_X1 _15942_ ( .A(\u_lsu.pmem[6214] ), .B1(_02325_ ), .B2(_02339_ ), .ZN(_02344_ ) );
BUF_X4 _15943_ ( .A(_10904_ ), .Z(_02345_ ) );
NAND4_X1 _15944_ ( .A1(_09957_ ), .A2(_11536_ ), .A3(_02313_ ), .A4(_02345_ ), .ZN(_02346_ ) );
AOI21_X1 _15945_ ( .A(fanout_net_29 ), .B1(_02344_ ), .B2(_02346_ ), .ZN(_00797_ ) );
OAI21_X1 _15946_ ( .A(\u_lsu.pmem[6213] ), .B1(_02325_ ), .B2(_02339_ ), .ZN(_02347_ ) );
BUF_X4 _15947_ ( .A(_11381_ ), .Z(_02348_ ) );
NAND4_X1 _15948_ ( .A1(_09961_ ), .A2(_11536_ ), .A3(_02348_ ), .A4(_02345_ ), .ZN(_02349_ ) );
AOI21_X1 _15949_ ( .A(fanout_net_29 ), .B1(_02347_ ), .B2(_02349_ ), .ZN(_00798_ ) );
OAI21_X1 _15950_ ( .A(\u_lsu.pmem[6212] ), .B1(_02325_ ), .B2(_02339_ ), .ZN(_02350_ ) );
NAND4_X1 _15951_ ( .A1(_09966_ ), .A2(_11536_ ), .A3(_02348_ ), .A4(_02345_ ), .ZN(_02351_ ) );
AOI21_X1 _15952_ ( .A(fanout_net_29 ), .B1(_02350_ ), .B2(_02351_ ), .ZN(_00799_ ) );
OAI21_X1 _15953_ ( .A(\u_lsu.pmem[6211] ), .B1(_02325_ ), .B2(_02339_ ), .ZN(_02352_ ) );
NAND4_X1 _15954_ ( .A1(_09970_ ), .A2(_11536_ ), .A3(_02348_ ), .A4(_02345_ ), .ZN(_02353_ ) );
AOI21_X1 _15955_ ( .A(fanout_net_29 ), .B1(_02352_ ), .B2(_02353_ ), .ZN(_00800_ ) );
OAI21_X1 _15956_ ( .A(\u_lsu.pmem[6210] ), .B1(_02325_ ), .B2(_02339_ ), .ZN(_02354_ ) );
NAND4_X1 _15957_ ( .A1(_09974_ ), .A2(_11536_ ), .A3(_02348_ ), .A4(_02345_ ), .ZN(_02355_ ) );
AOI21_X1 _15958_ ( .A(fanout_net_29 ), .B1(_02354_ ), .B2(_02355_ ), .ZN(_00801_ ) );
BUF_X4 _15959_ ( .A(_11582_ ), .Z(_02356_ ) );
OAI21_X1 _15960_ ( .A(\u_lsu.pmem[6209] ), .B1(_02356_ ), .B2(_02339_ ), .ZN(_02357_ ) );
NAND4_X1 _15961_ ( .A1(_09978_ ), .A2(_11536_ ), .A3(_02348_ ), .A4(_02345_ ), .ZN(_02358_ ) );
AOI21_X1 _15962_ ( .A(fanout_net_29 ), .B1(_02357_ ), .B2(_02358_ ), .ZN(_00802_ ) );
OAI21_X1 _15963_ ( .A(\u_lsu.pmem[6208] ), .B1(_02356_ ), .B2(_02339_ ), .ZN(_02359_ ) );
NAND4_X1 _15964_ ( .A1(_09982_ ), .A2(_11536_ ), .A3(_02348_ ), .A4(_02345_ ), .ZN(_02360_ ) );
AOI21_X1 _15965_ ( .A(fanout_net_29 ), .B1(_02359_ ), .B2(_02360_ ), .ZN(_00803_ ) );
NAND4_X1 _15966_ ( .A1(_09987_ ), .A2(_02286_ ), .A3(_02287_ ), .A4(_02279_ ), .ZN(_02361_ ) );
NAND3_X4 _15967_ ( .A1(_09135_ ), .A2(_09538_ ), .A3(_09989_ ), .ZN(_02362_ ) );
BUF_X4 _15968_ ( .A(_02362_ ), .Z(_02363_ ) );
OAI21_X1 _15969_ ( .A(\u_lsu.pmem[6183] ), .B1(_02277_ ), .B2(_02363_ ), .ZN(_02364_ ) );
AOI21_X1 _15970_ ( .A(fanout_net_29 ), .B1(_02361_ ), .B2(_02364_ ), .ZN(_00804_ ) );
NAND4_X1 _15971_ ( .A1(_09994_ ), .A2(_02286_ ), .A3(_02287_ ), .A4(_02279_ ), .ZN(_02365_ ) );
OAI21_X1 _15972_ ( .A(\u_lsu.pmem[6182] ), .B1(_02277_ ), .B2(_02363_ ), .ZN(_02366_ ) );
AOI21_X1 _15973_ ( .A(fanout_net_29 ), .B1(_02365_ ), .B2(_02366_ ), .ZN(_00805_ ) );
NAND4_X1 _15974_ ( .A1(_09997_ ), .A2(_02286_ ), .A3(_02287_ ), .A4(_02279_ ), .ZN(_02367_ ) );
OAI21_X1 _15975_ ( .A(\u_lsu.pmem[6181] ), .B1(_02277_ ), .B2(_02363_ ), .ZN(_02368_ ) );
AOI21_X1 _15976_ ( .A(fanout_net_29 ), .B1(_02367_ ), .B2(_02368_ ), .ZN(_00806_ ) );
NAND4_X1 _15977_ ( .A1(_09770_ ), .A2(_02286_ ), .A3(_09869_ ), .A4(_02279_ ), .ZN(_02369_ ) );
OAI21_X1 _15978_ ( .A(\u_lsu.pmem[4324] ), .B1(_02277_ ), .B2(_09751_ ), .ZN(_02370_ ) );
AOI21_X1 _15979_ ( .A(fanout_net_29 ), .B1(_02369_ ), .B2(_02370_ ), .ZN(_00807_ ) );
BUF_X4 _15980_ ( .A(_11492_ ), .Z(_02371_ ) );
NAND4_X1 _15981_ ( .A1(_10408_ ), .A2(_02225_ ), .A3(_02287_ ), .A4(_02371_ ), .ZN(_02372_ ) );
OAI21_X1 _15982_ ( .A(\u_lsu.pmem[3748] ), .B1(_02342_ ), .B2(_10399_ ), .ZN(_02373_ ) );
AOI21_X1 _15983_ ( .A(fanout_net_29 ), .B1(_02372_ ), .B2(_02373_ ), .ZN(_00808_ ) );
NOR2_X1 _15984_ ( .A1(_09641_ ), .A2(_02362_ ), .ZN(_02374_ ) );
OAI21_X1 _15985_ ( .A(_10715_ ), .B1(_02374_ ), .B2(\u_lsu.pmem[6180] ), .ZN(_02375_ ) );
AOI21_X1 _15986_ ( .A(_02375_ ), .B1(_09691_ ), .B2(_02374_ ), .ZN(_00809_ ) );
OAI21_X1 _15987_ ( .A(\u_lsu.pmem[6179] ), .B1(_02356_ ), .B2(_02363_ ), .ZN(_02376_ ) );
NAND4_X1 _15988_ ( .A1(_11385_ ), .A2(_02318_ ), .A3(_02348_ ), .A4(_10001_ ), .ZN(_02377_ ) );
AOI21_X1 _15989_ ( .A(fanout_net_29 ), .B1(_02376_ ), .B2(_02377_ ), .ZN(_00810_ ) );
OAI21_X1 _15990_ ( .A(\u_lsu.pmem[6178] ), .B1(_02356_ ), .B2(_02363_ ), .ZN(_02378_ ) );
BUF_X4 _15991_ ( .A(_09611_ ), .Z(_02379_ ) );
NAND4_X1 _15992_ ( .A1(_02379_ ), .A2(_02318_ ), .A3(_02348_ ), .A4(_10001_ ), .ZN(_02380_ ) );
AOI21_X1 _15993_ ( .A(fanout_net_29 ), .B1(_02378_ ), .B2(_02380_ ), .ZN(_00811_ ) );
OAI21_X1 _15994_ ( .A(\u_lsu.pmem[6177] ), .B1(_02356_ ), .B2(_02363_ ), .ZN(_02381_ ) );
BUF_X4 _15995_ ( .A(_10548_ ), .Z(_02382_ ) );
NAND4_X1 _15996_ ( .A1(_11414_ ), .A2(_02382_ ), .A3(_02348_ ), .A4(_10001_ ), .ZN(_02383_ ) );
AOI21_X1 _15997_ ( .A(fanout_net_29 ), .B1(_02381_ ), .B2(_02383_ ), .ZN(_00812_ ) );
NAND4_X1 _15998_ ( .A1(_10021_ ), .A2(_02286_ ), .A3(_02287_ ), .A4(_02279_ ), .ZN(_02384_ ) );
BUF_X4 _15999_ ( .A(_02209_ ), .Z(_02385_ ) );
OAI21_X1 _16000_ ( .A(\u_lsu.pmem[6176] ), .B1(_02385_ ), .B2(_02363_ ), .ZN(_02386_ ) );
AOI21_X1 _16001_ ( .A(fanout_net_29 ), .B1(_02384_ ), .B2(_02386_ ), .ZN(_00813_ ) );
BUF_X4 _16002_ ( .A(_09133_ ), .Z(_02387_ ) );
NAND4_X1 _16003_ ( .A1(_02387_ ), .A2(_11423_ ), .A3(_10824_ ), .A4(\alu_result_out[8] ), .ZN(_02388_ ) );
NAND3_X1 _16004_ ( .A1(_09116_ ), .A2(_09805_ ), .A3(_09605_ ), .ZN(_02389_ ) );
BUF_X4 _16005_ ( .A(_02389_ ), .Z(_02390_ ) );
OAI21_X1 _16006_ ( .A(\u_lsu.pmem[6151] ), .B1(_02390_ ), .B2(_11019_ ), .ZN(_02391_ ) );
AOI21_X1 _16007_ ( .A(fanout_net_29 ), .B1(_02388_ ), .B2(_02391_ ), .ZN(_00814_ ) );
NAND4_X1 _16008_ ( .A1(_02387_ ), .A2(_10444_ ), .A3(_10824_ ), .A4(\alu_result_out[8] ), .ZN(_02392_ ) );
OAI21_X1 _16009_ ( .A(\u_lsu.pmem[6150] ), .B1(_02390_ ), .B2(_11019_ ), .ZN(_02393_ ) );
AOI21_X1 _16010_ ( .A(fanout_net_29 ), .B1(_02392_ ), .B2(_02393_ ), .ZN(_00815_ ) );
NAND4_X1 _16011_ ( .A1(_02387_ ), .A2(_10448_ ), .A3(_10824_ ), .A4(\alu_result_out[8] ), .ZN(_02394_ ) );
OAI21_X1 _16012_ ( .A(\u_lsu.pmem[6149] ), .B1(_02390_ ), .B2(_11019_ ), .ZN(_02395_ ) );
AOI21_X1 _16013_ ( .A(fanout_net_29 ), .B1(_02394_ ), .B2(_02395_ ), .ZN(_00816_ ) );
NOR2_X1 _16014_ ( .A1(_02389_ ), .A2(_10012_ ), .ZN(_02396_ ) );
NOR2_X1 _16015_ ( .A1(_02396_ ), .A2(\u_lsu.pmem[6148] ), .ZN(_02397_ ) );
AOI211_X1 _16016_ ( .A(fanout_net_29 ), .B(_02397_ ), .C1(_09146_ ), .C2(_02396_ ), .ZN(_00817_ ) );
NAND4_X1 _16017_ ( .A1(_02387_ ), .A2(_10456_ ), .A3(_10824_ ), .A4(\alu_result_out[8] ), .ZN(_02398_ ) );
OAI21_X1 _16018_ ( .A(\u_lsu.pmem[6147] ), .B1(_02390_ ), .B2(_11019_ ), .ZN(_02399_ ) );
AOI21_X1 _16019_ ( .A(fanout_net_29 ), .B1(_02398_ ), .B2(_02399_ ), .ZN(_00818_ ) );
NAND4_X1 _16020_ ( .A1(_10411_ ), .A2(_02225_ ), .A3(_02287_ ), .A4(_02371_ ), .ZN(_02400_ ) );
OAI21_X1 _16021_ ( .A(\u_lsu.pmem[3747] ), .B1(_02342_ ), .B2(_10399_ ), .ZN(_02401_ ) );
AOI21_X1 _16022_ ( .A(fanout_net_29 ), .B1(_02400_ ), .B2(_02401_ ), .ZN(_00819_ ) );
BUF_X4 _16023_ ( .A(_09673_ ), .Z(_02402_ ) );
NAND4_X1 _16024_ ( .A1(_11021_ ), .A2(_02225_ ), .A3(_02402_ ), .A4(_02279_ ), .ZN(_02403_ ) );
OAI21_X1 _16025_ ( .A(\u_lsu.pmem[6146] ), .B1(_02390_ ), .B2(_11019_ ), .ZN(_02404_ ) );
AOI21_X1 _16026_ ( .A(fanout_net_30 ), .B1(_02403_ ), .B2(_02404_ ), .ZN(_00820_ ) );
NAND4_X1 _16027_ ( .A1(_02387_ ), .A2(_10463_ ), .A3(_10824_ ), .A4(_09607_ ), .ZN(_02405_ ) );
OAI21_X1 _16028_ ( .A(\u_lsu.pmem[6145] ), .B1(_02390_ ), .B2(_11019_ ), .ZN(_02406_ ) );
AOI21_X1 _16029_ ( .A(fanout_net_30 ), .B1(_02405_ ), .B2(_02406_ ), .ZN(_00821_ ) );
NAND4_X1 _16030_ ( .A1(_02387_ ), .A2(_10467_ ), .A3(_10824_ ), .A4(_09607_ ), .ZN(_02407_ ) );
OAI21_X1 _16031_ ( .A(\u_lsu.pmem[6144] ), .B1(_02390_ ), .B2(_09496_ ), .ZN(_02408_ ) );
AOI21_X1 _16032_ ( .A(fanout_net_30 ), .B1(_02407_ ), .B2(_02408_ ), .ZN(_00822_ ) );
BUF_X2 _16033_ ( .A(_09020_ ), .Z(_02409_ ) );
NAND3_X1 _16034_ ( .A1(_10054_ ), .A2(_02409_ ), .A3(_10055_ ), .ZN(_02410_ ) );
BUF_X4 _16035_ ( .A(_02410_ ), .Z(_02411_ ) );
OAI21_X1 _16036_ ( .A(\u_lsu.pmem[6119] ), .B1(_02356_ ), .B2(_02411_ ), .ZN(_02412_ ) );
CLKBUF_X2 _16037_ ( .A(_09493_ ), .Z(_02413_ ) );
OR4_X1 _16038_ ( .A1(_09565_ ), .A2(_09499_ ), .A3(_02413_ ), .A4(_02410_ ), .ZN(_02414_ ) );
AOI21_X1 _16039_ ( .A(fanout_net_30 ), .B1(_02412_ ), .B2(_02414_ ), .ZN(_00823_ ) );
BUF_X4 _16040_ ( .A(_11334_ ), .Z(_02415_ ) );
NAND4_X1 _16041_ ( .A1(_10062_ ), .A2(_02225_ ), .A3(_02402_ ), .A4(_02415_ ), .ZN(_02416_ ) );
OAI21_X1 _16042_ ( .A(\u_lsu.pmem[6118] ), .B1(_02385_ ), .B2(_02411_ ), .ZN(_02417_ ) );
AOI21_X1 _16043_ ( .A(fanout_net_30 ), .B1(_02416_ ), .B2(_02417_ ), .ZN(_00824_ ) );
NAND4_X1 _16044_ ( .A1(_10075_ ), .A2(_02225_ ), .A3(_02402_ ), .A4(_02415_ ), .ZN(_02418_ ) );
OAI21_X1 _16045_ ( .A(\u_lsu.pmem[6117] ), .B1(_02385_ ), .B2(_02411_ ), .ZN(_02419_ ) );
AOI21_X1 _16046_ ( .A(fanout_net_30 ), .B1(_02418_ ), .B2(_02419_ ), .ZN(_00825_ ) );
BUF_X4 _16047_ ( .A(_10886_ ), .Z(_02420_ ) );
NAND4_X1 _16048_ ( .A1(_10079_ ), .A2(_02420_ ), .A3(_02402_ ), .A4(_02415_ ), .ZN(_02421_ ) );
OAI21_X1 _16049_ ( .A(\u_lsu.pmem[6116] ), .B1(_02385_ ), .B2(_02411_ ), .ZN(_02422_ ) );
AOI21_X1 _16050_ ( .A(fanout_net_30 ), .B1(_02421_ ), .B2(_02422_ ), .ZN(_00826_ ) );
NAND4_X1 _16051_ ( .A1(_10084_ ), .A2(_02420_ ), .A3(_02402_ ), .A4(_02415_ ), .ZN(_02423_ ) );
OAI21_X1 _16052_ ( .A(\u_lsu.pmem[6115] ), .B1(_02385_ ), .B2(_02411_ ), .ZN(_02424_ ) );
AOI21_X1 _16053_ ( .A(fanout_net_30 ), .B1(_02423_ ), .B2(_02424_ ), .ZN(_00827_ ) );
NAND4_X1 _16054_ ( .A1(_10088_ ), .A2(_02420_ ), .A3(_02402_ ), .A4(_02415_ ), .ZN(_02425_ ) );
OAI21_X1 _16055_ ( .A(\u_lsu.pmem[6114] ), .B1(_02385_ ), .B2(_02411_ ), .ZN(_02426_ ) );
AOI21_X1 _16056_ ( .A(fanout_net_30 ), .B1(_02425_ ), .B2(_02426_ ), .ZN(_00828_ ) );
NAND4_X1 _16057_ ( .A1(_10094_ ), .A2(_02420_ ), .A3(_02402_ ), .A4(_02415_ ), .ZN(_02427_ ) );
OAI21_X1 _16058_ ( .A(\u_lsu.pmem[6113] ), .B1(_02385_ ), .B2(_02411_ ), .ZN(_02428_ ) );
AOI21_X1 _16059_ ( .A(fanout_net_30 ), .B1(_02427_ ), .B2(_02428_ ), .ZN(_00829_ ) );
BUF_X4 _16060_ ( .A(_02196_ ), .Z(_02429_ ) );
NAND4_X1 _16061_ ( .A1(_10414_ ), .A2(_02420_ ), .A3(_02429_ ), .A4(_02371_ ), .ZN(_02430_ ) );
OAI21_X1 _16062_ ( .A(\u_lsu.pmem[3746] ), .B1(_02342_ ), .B2(_10399_ ), .ZN(_02431_ ) );
AOI21_X1 _16063_ ( .A(fanout_net_30 ), .B1(_02430_ ), .B2(_02431_ ), .ZN(_00830_ ) );
NAND4_X1 _16064_ ( .A1(_10098_ ), .A2(_02420_ ), .A3(_02402_ ), .A4(_02415_ ), .ZN(_02432_ ) );
OAI21_X1 _16065_ ( .A(\u_lsu.pmem[6112] ), .B1(_02385_ ), .B2(_02411_ ), .ZN(_02433_ ) );
AOI21_X1 _16066_ ( .A(fanout_net_30 ), .B1(_02432_ ), .B2(_02433_ ), .ZN(_00831_ ) );
NAND3_X1 _16067_ ( .A1(_10103_ ), .A2(_02409_ ), .A3(_10055_ ), .ZN(_02434_ ) );
BUF_X4 _16068_ ( .A(_02434_ ), .Z(_02435_ ) );
OAI21_X1 _16069_ ( .A(\u_lsu.pmem[6087] ), .B1(_02356_ ), .B2(_02435_ ), .ZN(_02436_ ) );
OR4_X1 _16070_ ( .A1(_09565_ ), .A2(_09499_ ), .A3(_02413_ ), .A4(_02434_ ), .ZN(_02437_ ) );
AOI21_X1 _16071_ ( .A(fanout_net_30 ), .B1(_02436_ ), .B2(_02437_ ), .ZN(_00832_ ) );
NAND4_X1 _16072_ ( .A1(_10117_ ), .A2(_02420_ ), .A3(_02402_ ), .A4(_02415_ ), .ZN(_02438_ ) );
OAI21_X1 _16073_ ( .A(\u_lsu.pmem[6086] ), .B1(_02385_ ), .B2(_02435_ ), .ZN(_02439_ ) );
AOI21_X1 _16074_ ( .A(fanout_net_30 ), .B1(_02438_ ), .B2(_02439_ ), .ZN(_00833_ ) );
NAND4_X1 _16075_ ( .A1(_10121_ ), .A2(_02420_ ), .A3(_02402_ ), .A4(_02415_ ), .ZN(_02440_ ) );
OAI21_X1 _16076_ ( .A(\u_lsu.pmem[6085] ), .B1(_02385_ ), .B2(_02435_ ), .ZN(_02441_ ) );
AOI21_X1 _16077_ ( .A(fanout_net_30 ), .B1(_02440_ ), .B2(_02441_ ), .ZN(_00834_ ) );
BUF_X4 _16078_ ( .A(_09673_ ), .Z(_02442_ ) );
NAND4_X1 _16079_ ( .A1(_10125_ ), .A2(_02420_ ), .A3(_02442_ ), .A4(_02415_ ), .ZN(_02443_ ) );
BUF_X4 _16080_ ( .A(_02209_ ), .Z(_02444_ ) );
OAI21_X1 _16081_ ( .A(\u_lsu.pmem[6084] ), .B1(_02444_ ), .B2(_02435_ ), .ZN(_02445_ ) );
AOI21_X1 _16082_ ( .A(fanout_net_30 ), .B1(_02443_ ), .B2(_02445_ ), .ZN(_00835_ ) );
BUF_X4 _16083_ ( .A(_11334_ ), .Z(_02446_ ) );
NAND4_X1 _16084_ ( .A1(_10131_ ), .A2(_02420_ ), .A3(_02442_ ), .A4(_02446_ ), .ZN(_02447_ ) );
OAI21_X1 _16085_ ( .A(\u_lsu.pmem[6083] ), .B1(_02444_ ), .B2(_02435_ ), .ZN(_02448_ ) );
AOI21_X1 _16086_ ( .A(fanout_net_30 ), .B1(_02447_ ), .B2(_02448_ ), .ZN(_00836_ ) );
BUF_X4 _16087_ ( .A(_10886_ ), .Z(_02449_ ) );
NAND4_X1 _16088_ ( .A1(_10135_ ), .A2(_02449_ ), .A3(_02442_ ), .A4(_02446_ ), .ZN(_02450_ ) );
OAI21_X1 _16089_ ( .A(\u_lsu.pmem[6082] ), .B1(_02444_ ), .B2(_02435_ ), .ZN(_02451_ ) );
AOI21_X1 _16090_ ( .A(fanout_net_30 ), .B1(_02450_ ), .B2(_02451_ ), .ZN(_00837_ ) );
NAND4_X1 _16091_ ( .A1(_10138_ ), .A2(_02449_ ), .A3(_02442_ ), .A4(_02446_ ), .ZN(_02452_ ) );
OAI21_X1 _16092_ ( .A(\u_lsu.pmem[6081] ), .B1(_02444_ ), .B2(_02435_ ), .ZN(_02453_ ) );
AOI21_X1 _16093_ ( .A(fanout_net_30 ), .B1(_02452_ ), .B2(_02453_ ), .ZN(_00838_ ) );
NAND4_X1 _16094_ ( .A1(_10144_ ), .A2(_02449_ ), .A3(_02442_ ), .A4(_02446_ ), .ZN(_02454_ ) );
OAI21_X1 _16095_ ( .A(\u_lsu.pmem[6080] ), .B1(_02444_ ), .B2(_02435_ ), .ZN(_02455_ ) );
AOI21_X1 _16096_ ( .A(fanout_net_30 ), .B1(_02454_ ), .B2(_02455_ ), .ZN(_00839_ ) );
NAND4_X1 _16097_ ( .A1(_10148_ ), .A2(_02449_ ), .A3(_02442_ ), .A4(_02446_ ), .ZN(_02456_ ) );
BUF_X4 _16098_ ( .A(_09020_ ), .Z(_02457_ ) );
AND3_X1 _16099_ ( .A1(_09488_ ), .A2(_02457_ ), .A3(_10055_ ), .ZN(_02458_ ) );
INV_X1 _16100_ ( .A(_02458_ ), .ZN(_02459_ ) );
BUF_X4 _16101_ ( .A(_02459_ ), .Z(_02460_ ) );
OAI21_X1 _16102_ ( .A(\u_lsu.pmem[6055] ), .B1(_02444_ ), .B2(_02460_ ), .ZN(_02461_ ) );
AOI21_X1 _16103_ ( .A(fanout_net_30 ), .B1(_02456_ ), .B2(_02461_ ), .ZN(_00840_ ) );
NAND4_X1 _16104_ ( .A1(_10417_ ), .A2(_02449_ ), .A3(_02429_ ), .A4(_02371_ ), .ZN(_02462_ ) );
OAI21_X1 _16105_ ( .A(\u_lsu.pmem[3745] ), .B1(_02342_ ), .B2(_10399_ ), .ZN(_02463_ ) );
AOI21_X1 _16106_ ( .A(fanout_net_30 ), .B1(_02462_ ), .B2(_02463_ ), .ZN(_00841_ ) );
NAND4_X1 _16107_ ( .A1(_10156_ ), .A2(_02449_ ), .A3(_02442_ ), .A4(_02446_ ), .ZN(_02464_ ) );
OAI21_X1 _16108_ ( .A(\u_lsu.pmem[6054] ), .B1(_02444_ ), .B2(_02460_ ), .ZN(_02465_ ) );
AOI21_X1 _16109_ ( .A(fanout_net_30 ), .B1(_02464_ ), .B2(_02465_ ), .ZN(_00842_ ) );
NAND4_X1 _16110_ ( .A1(_10160_ ), .A2(_02449_ ), .A3(_02442_ ), .A4(_02446_ ), .ZN(_02466_ ) );
OAI21_X1 _16111_ ( .A(\u_lsu.pmem[6053] ), .B1(_02444_ ), .B2(_02460_ ), .ZN(_02467_ ) );
AOI21_X1 _16112_ ( .A(fanout_net_30 ), .B1(_02466_ ), .B2(_02467_ ), .ZN(_00843_ ) );
NAND4_X1 _16113_ ( .A1(_10166_ ), .A2(_02449_ ), .A3(_02442_ ), .A4(_02446_ ), .ZN(_02468_ ) );
OAI21_X1 _16114_ ( .A(\u_lsu.pmem[6052] ), .B1(_02444_ ), .B2(_02460_ ), .ZN(_02469_ ) );
AOI21_X1 _16115_ ( .A(fanout_net_30 ), .B1(_02468_ ), .B2(_02469_ ), .ZN(_00844_ ) );
NAND4_X1 _16116_ ( .A1(_10169_ ), .A2(_02449_ ), .A3(_02442_ ), .A4(_02446_ ), .ZN(_02470_ ) );
OAI21_X1 _16117_ ( .A(\u_lsu.pmem[6051] ), .B1(_02444_ ), .B2(_02460_ ), .ZN(_02471_ ) );
AOI21_X1 _16118_ ( .A(fanout_net_30 ), .B1(_02470_ ), .B2(_02471_ ), .ZN(_00845_ ) );
BUF_X4 _16119_ ( .A(_09673_ ), .Z(_02472_ ) );
NAND4_X1 _16120_ ( .A1(_10172_ ), .A2(_02449_ ), .A3(_02472_ ), .A4(_02446_ ), .ZN(_02473_ ) );
BUF_X4 _16121_ ( .A(_02209_ ), .Z(_02474_ ) );
OAI21_X1 _16122_ ( .A(\u_lsu.pmem[6050] ), .B1(_02474_ ), .B2(_02460_ ), .ZN(_02475_ ) );
AOI21_X1 _16123_ ( .A(fanout_net_30 ), .B1(_02473_ ), .B2(_02475_ ), .ZN(_00846_ ) );
BUF_X4 _16124_ ( .A(_10886_ ), .Z(_02476_ ) );
BUF_X4 _16125_ ( .A(_11334_ ), .Z(_02477_ ) );
NAND4_X1 _16126_ ( .A1(_10176_ ), .A2(_02476_ ), .A3(_02472_ ), .A4(_02477_ ), .ZN(_02478_ ) );
OAI21_X1 _16127_ ( .A(\u_lsu.pmem[6049] ), .B1(_02474_ ), .B2(_02460_ ), .ZN(_02479_ ) );
AOI21_X1 _16128_ ( .A(fanout_net_30 ), .B1(_02478_ ), .B2(_02479_ ), .ZN(_00847_ ) );
OAI21_X1 _16129_ ( .A(\u_lsu.pmem[6048] ), .B1(_02356_ ), .B2(_02460_ ), .ZN(_02480_ ) );
CLKBUF_X2 _16130_ ( .A(_09493_ ), .Z(_02481_ ) );
OR4_X1 _16131_ ( .A1(_09497_ ), .A2(_02459_ ), .A3(_09498_ ), .A4(_02481_ ), .ZN(_02482_ ) );
AOI21_X1 _16132_ ( .A(fanout_net_30 ), .B1(_02480_ ), .B2(_02482_ ), .ZN(_00848_ ) );
BUF_X4 _16133_ ( .A(_09601_ ), .Z(_02483_ ) );
BUF_X4 _16134_ ( .A(_02457_ ), .Z(_02484_ ) );
BUF_X4 _16135_ ( .A(_02484_ ), .Z(_02485_ ) );
BUF_X4 _16136_ ( .A(_02485_ ), .Z(_02486_ ) );
NAND4_X1 _16137_ ( .A1(_02483_ ), .A2(_11423_ ), .A3(_02486_ ), .A4(_02477_ ), .ZN(_02487_ ) );
NAND3_X1 _16138_ ( .A1(_09595_ ), .A2(_02484_ ), .A3(_09875_ ), .ZN(_02488_ ) );
BUF_X4 _16139_ ( .A(_02488_ ), .Z(_02489_ ) );
OAI21_X1 _16140_ ( .A(\u_lsu.pmem[6023] ), .B1(_02489_ ), .B2(_11337_ ), .ZN(_02490_ ) );
AOI21_X1 _16141_ ( .A(fanout_net_30 ), .B1(_02487_ ), .B2(_02490_ ), .ZN(_00849_ ) );
NAND4_X1 _16142_ ( .A1(_02483_ ), .A2(_10444_ ), .A3(_02486_ ), .A4(_02477_ ), .ZN(_02491_ ) );
BUF_X4 _16143_ ( .A(_09515_ ), .Z(_02492_ ) );
OAI21_X1 _16144_ ( .A(\u_lsu.pmem[6022] ), .B1(_02489_ ), .B2(_02492_ ), .ZN(_02493_ ) );
AOI21_X1 _16145_ ( .A(fanout_net_31 ), .B1(_02491_ ), .B2(_02493_ ), .ZN(_00850_ ) );
NAND4_X1 _16146_ ( .A1(_02483_ ), .A2(_10448_ ), .A3(_02486_ ), .A4(_02477_ ), .ZN(_02494_ ) );
OAI21_X1 _16147_ ( .A(\u_lsu.pmem[6021] ), .B1(_02489_ ), .B2(_02492_ ), .ZN(_02495_ ) );
AOI21_X1 _16148_ ( .A(fanout_net_31 ), .B1(_02494_ ), .B2(_02495_ ), .ZN(_00851_ ) );
NAND4_X1 _16149_ ( .A1(_10018_ ), .A2(_11212_ ), .A3(_09944_ ), .A4(_10398_ ), .ZN(_02496_ ) );
OAI21_X1 _16150_ ( .A(\u_lsu.pmem[3744] ), .B1(_02342_ ), .B2(_10399_ ), .ZN(_02497_ ) );
AOI21_X1 _16151_ ( .A(fanout_net_31 ), .B1(_02496_ ), .B2(_02497_ ), .ZN(_00852_ ) );
NAND4_X1 _16152_ ( .A1(_02483_ ), .A2(_10453_ ), .A3(_02486_ ), .A4(_02477_ ), .ZN(_02498_ ) );
OAI21_X1 _16153_ ( .A(\u_lsu.pmem[6020] ), .B1(_02489_ ), .B2(_02492_ ), .ZN(_02499_ ) );
AOI21_X1 _16154_ ( .A(fanout_net_31 ), .B1(_02498_ ), .B2(_02499_ ), .ZN(_00853_ ) );
BUF_X4 _16155_ ( .A(_02485_ ), .Z(_02500_ ) );
NAND4_X1 _16156_ ( .A1(_02483_ ), .A2(_10456_ ), .A3(_02500_ ), .A4(_02477_ ), .ZN(_02501_ ) );
OAI21_X1 _16157_ ( .A(\u_lsu.pmem[6019] ), .B1(_02489_ ), .B2(_02492_ ), .ZN(_02502_ ) );
AOI21_X1 _16158_ ( .A(fanout_net_31 ), .B1(_02501_ ), .B2(_02502_ ), .ZN(_00854_ ) );
OAI21_X1 _16159_ ( .A(\u_lsu.pmem[6018] ), .B1(_02489_ ), .B2(_02189_ ), .ZN(_02503_ ) );
NAND4_X1 _16160_ ( .A1(_09874_ ), .A2(_10976_ ), .A3(_09909_ ), .A4(_02345_ ), .ZN(_02504_ ) );
AOI21_X1 _16161_ ( .A(fanout_net_31 ), .B1(_02503_ ), .B2(_02504_ ), .ZN(_00855_ ) );
NAND4_X1 _16162_ ( .A1(_02483_ ), .A2(_10463_ ), .A3(_02500_ ), .A4(_02477_ ), .ZN(_02505_ ) );
OAI21_X1 _16163_ ( .A(\u_lsu.pmem[6017] ), .B1(_02489_ ), .B2(_02492_ ), .ZN(_02506_ ) );
AOI21_X1 _16164_ ( .A(fanout_net_31 ), .B1(_02505_ ), .B2(_02506_ ), .ZN(_00856_ ) );
NAND4_X1 _16165_ ( .A1(_02483_ ), .A2(_10467_ ), .A3(_02500_ ), .A4(_02477_ ), .ZN(_02507_ ) );
OAI21_X1 _16166_ ( .A(\u_lsu.pmem[6016] ), .B1(_02489_ ), .B2(_02492_ ), .ZN(_02508_ ) );
AOI21_X1 _16167_ ( .A(fanout_net_31 ), .B1(_02507_ ), .B2(_02508_ ), .ZN(_00857_ ) );
AND3_X2 _16168_ ( .A1(_10008_ ), .A2(_09020_ ), .A3(_10009_ ), .ZN(_02509_ ) );
INV_X1 _16169_ ( .A(_02509_ ), .ZN(_02510_ ) );
BUF_X4 _16170_ ( .A(_02510_ ), .Z(_02511_ ) );
BUF_X4 _16171_ ( .A(_02511_ ), .Z(_02512_ ) );
OAI21_X1 _16172_ ( .A(\u_lsu.pmem[5991] ), .B1(_02356_ ), .B2(_02512_ ), .ZN(_02513_ ) );
OR4_X1 _16173_ ( .A1(_09565_ ), .A2(_09499_ ), .A3(_02413_ ), .A4(_02511_ ), .ZN(_02514_ ) );
AOI21_X1 _16174_ ( .A(fanout_net_31 ), .B1(_02513_ ), .B2(_02514_ ), .ZN(_00858_ ) );
OAI21_X1 _16175_ ( .A(\u_lsu.pmem[5990] ), .B1(_02356_ ), .B2(_02512_ ), .ZN(_02515_ ) );
OR4_X1 _16176_ ( .A1(_09576_ ), .A2(_09499_ ), .A3(_02413_ ), .A4(_02511_ ), .ZN(_02516_ ) );
AOI21_X1 _16177_ ( .A(fanout_net_31 ), .B1(_02515_ ), .B2(_02516_ ), .ZN(_00859_ ) );
BUF_X4 _16178_ ( .A(_11582_ ), .Z(_02517_ ) );
OAI21_X1 _16179_ ( .A(\u_lsu.pmem[5989] ), .B1(_02517_ ), .B2(_02512_ ), .ZN(_02518_ ) );
OR4_X1 _16180_ ( .A1(_09583_ ), .A2(_09499_ ), .A3(_02413_ ), .A4(_02511_ ), .ZN(_02519_ ) );
AOI21_X1 _16181_ ( .A(fanout_net_31 ), .B1(_02518_ ), .B2(_02519_ ), .ZN(_00860_ ) );
OAI21_X1 _16182_ ( .A(\u_lsu.pmem[5988] ), .B1(_02517_ ), .B2(_02512_ ), .ZN(_02520_ ) );
OR4_X1 _16183_ ( .A1(_09146_ ), .A2(_09499_ ), .A3(_02413_ ), .A4(_02510_ ), .ZN(_02521_ ) );
AOI21_X1 _16184_ ( .A(fanout_net_31 ), .B1(_02520_ ), .B2(_02521_ ), .ZN(_00861_ ) );
OAI21_X1 _16185_ ( .A(\u_lsu.pmem[5987] ), .B1(_02517_ ), .B2(_02512_ ), .ZN(_02522_ ) );
CLKBUF_X2 _16186_ ( .A(_09493_ ), .Z(_02523_ ) );
OR4_X1 _16187_ ( .A1(_09969_ ), .A2(_09499_ ), .A3(_02523_ ), .A4(_02510_ ), .ZN(_02524_ ) );
AOI21_X1 _16188_ ( .A(fanout_net_31 ), .B1(_02522_ ), .B2(_02524_ ), .ZN(_00862_ ) );
OAI21_X1 _16189_ ( .A(\u_lsu.pmem[3719] ), .B1(_10426_ ), .B2(_09911_ ), .ZN(_02525_ ) );
BUF_X4 _16190_ ( .A(_09522_ ), .Z(_02526_ ) );
NAND4_X1 _16191_ ( .A1(_10436_ ), .A2(_10976_ ), .A3(_02348_ ), .A4(_02526_ ), .ZN(_02527_ ) );
AOI21_X1 _16192_ ( .A(fanout_net_31 ), .B1(_02525_ ), .B2(_02527_ ), .ZN(_00863_ ) );
OAI21_X1 _16193_ ( .A(\u_lsu.pmem[5986] ), .B1(_02517_ ), .B2(_02512_ ), .ZN(_02528_ ) );
OR4_X1 _16194_ ( .A1(_09973_ ), .A2(_09499_ ), .A3(_02523_ ), .A4(_02510_ ), .ZN(_02529_ ) );
AOI21_X1 _16195_ ( .A(fanout_net_31 ), .B1(_02528_ ), .B2(_02529_ ), .ZN(_00864_ ) );
OAI21_X1 _16196_ ( .A(\u_lsu.pmem[5985] ), .B1(_02517_ ), .B2(_02512_ ), .ZN(_02530_ ) );
CLKBUF_X2 _16197_ ( .A(_09498_ ), .Z(_02531_ ) );
OR4_X1 _16198_ ( .A1(_09977_ ), .A2(_02531_ ), .A3(_02523_ ), .A4(_02510_ ), .ZN(_02532_ ) );
AOI21_X1 _16199_ ( .A(fanout_net_31 ), .B1(_02530_ ), .B2(_02532_ ), .ZN(_00865_ ) );
OAI21_X1 _16200_ ( .A(\u_lsu.pmem[5984] ), .B1(_02517_ ), .B2(_02512_ ), .ZN(_02533_ ) );
OR4_X1 _16201_ ( .A1(_09497_ ), .A2(_02531_ ), .A3(_02523_ ), .A4(_02510_ ), .ZN(_02534_ ) );
AOI21_X1 _16202_ ( .A(fanout_net_31 ), .B1(_02533_ ), .B2(_02534_ ), .ZN(_00866_ ) );
AND3_X2 _16203_ ( .A1(_10226_ ), .A2(_09020_ ), .A3(_10009_ ), .ZN(_02535_ ) );
INV_X1 _16204_ ( .A(_02535_ ), .ZN(_02536_ ) );
BUF_X4 _16205_ ( .A(_02536_ ), .Z(_02537_ ) );
BUF_X4 _16206_ ( .A(_02537_ ), .Z(_02538_ ) );
OAI21_X1 _16207_ ( .A(\u_lsu.pmem[5959] ), .B1(_02517_ ), .B2(_02538_ ), .ZN(_02539_ ) );
OR4_X1 _16208_ ( .A1(_09565_ ), .A2(_02531_ ), .A3(_02523_ ), .A4(_02537_ ), .ZN(_02540_ ) );
AOI21_X1 _16209_ ( .A(fanout_net_31 ), .B1(_02539_ ), .B2(_02540_ ), .ZN(_00867_ ) );
OAI21_X1 _16210_ ( .A(\u_lsu.pmem[5958] ), .B1(_02517_ ), .B2(_02538_ ), .ZN(_02541_ ) );
OR4_X1 _16211_ ( .A1(_09576_ ), .A2(_02531_ ), .A3(_02523_ ), .A4(_02537_ ), .ZN(_02542_ ) );
AOI21_X1 _16212_ ( .A(fanout_net_31 ), .B1(_02541_ ), .B2(_02542_ ), .ZN(_00868_ ) );
OAI21_X1 _16213_ ( .A(\u_lsu.pmem[5957] ), .B1(_02517_ ), .B2(_02538_ ), .ZN(_02543_ ) );
OR4_X1 _16214_ ( .A1(_09583_ ), .A2(_02531_ ), .A3(_02523_ ), .A4(_02537_ ), .ZN(_02544_ ) );
AOI21_X1 _16215_ ( .A(fanout_net_31 ), .B1(_02543_ ), .B2(_02544_ ), .ZN(_00869_ ) );
OAI21_X1 _16216_ ( .A(\u_lsu.pmem[5956] ), .B1(_02517_ ), .B2(_02538_ ), .ZN(_02545_ ) );
OR4_X1 _16217_ ( .A1(_09146_ ), .A2(_02531_ ), .A3(_02523_ ), .A4(_02536_ ), .ZN(_02546_ ) );
AOI21_X1 _16218_ ( .A(fanout_net_31 ), .B1(_02545_ ), .B2(_02546_ ), .ZN(_00870_ ) );
BUF_X4 _16219_ ( .A(_11582_ ), .Z(_02547_ ) );
OAI21_X1 _16220_ ( .A(\u_lsu.pmem[5955] ), .B1(_02547_ ), .B2(_02538_ ), .ZN(_02548_ ) );
OR4_X1 _16221_ ( .A1(_09969_ ), .A2(_02531_ ), .A3(_02523_ ), .A4(_02536_ ), .ZN(_02549_ ) );
AOI21_X1 _16222_ ( .A(fanout_net_31 ), .B1(_02548_ ), .B2(_02549_ ), .ZN(_00871_ ) );
OAI21_X1 _16223_ ( .A(\u_lsu.pmem[5954] ), .B1(_02547_ ), .B2(_02538_ ), .ZN(_02550_ ) );
OR4_X1 _16224_ ( .A1(_09973_ ), .A2(_02531_ ), .A3(_02523_ ), .A4(_02536_ ), .ZN(_02551_ ) );
AOI21_X1 _16225_ ( .A(fanout_net_31 ), .B1(_02550_ ), .B2(_02551_ ), .ZN(_00872_ ) );
OAI21_X1 _16226_ ( .A(\u_lsu.pmem[5953] ), .B1(_02547_ ), .B2(_02538_ ), .ZN(_02552_ ) );
OR4_X1 _16227_ ( .A1(_09977_ ), .A2(_02531_ ), .A3(_02481_ ), .A4(_02536_ ), .ZN(_02553_ ) );
AOI21_X1 _16228_ ( .A(fanout_net_31 ), .B1(_02552_ ), .B2(_02553_ ), .ZN(_00873_ ) );
NAND4_X1 _16229_ ( .A1(_10443_ ), .A2(_09658_ ), .A3(_02429_ ), .A4(_02371_ ), .ZN(_02554_ ) );
OAI21_X1 _16230_ ( .A(\u_lsu.pmem[3718] ), .B1(_10425_ ), .B2(_09984_ ), .ZN(_02555_ ) );
AOI21_X1 _16231_ ( .A(fanout_net_31 ), .B1(_02554_ ), .B2(_02555_ ), .ZN(_00874_ ) );
OAI21_X1 _16232_ ( .A(\u_lsu.pmem[5952] ), .B1(_02547_ ), .B2(_02538_ ), .ZN(_02556_ ) );
OR4_X1 _16233_ ( .A1(_09497_ ), .A2(_02531_ ), .A3(_02481_ ), .A4(_02536_ ), .ZN(_02557_ ) );
AOI21_X1 _16234_ ( .A(fanout_net_31 ), .B1(_02556_ ), .B2(_02557_ ), .ZN(_00875_ ) );
NAND4_X1 _16235_ ( .A1(_10250_ ), .A2(_02476_ ), .A3(_02472_ ), .A4(_02477_ ), .ZN(_02558_ ) );
AND3_X1 _16236_ ( .A1(_10253_ ), .A2(_09020_ ), .A3(_10744_ ), .ZN(_02559_ ) );
INV_X1 _16237_ ( .A(_02559_ ), .ZN(_02560_ ) );
BUF_X4 _16238_ ( .A(_02560_ ), .Z(_02561_ ) );
OAI21_X1 _16239_ ( .A(\u_lsu.pmem[5927] ), .B1(_02474_ ), .B2(_02561_ ), .ZN(_02562_ ) );
AOI21_X1 _16240_ ( .A(fanout_net_31 ), .B1(_02558_ ), .B2(_02562_ ), .ZN(_00876_ ) );
NAND4_X1 _16241_ ( .A1(_10263_ ), .A2(_02476_ ), .A3(_02472_ ), .A4(_02477_ ), .ZN(_02563_ ) );
OAI21_X1 _16242_ ( .A(\u_lsu.pmem[5926] ), .B1(_02474_ ), .B2(_02561_ ), .ZN(_02564_ ) );
AOI21_X1 _16243_ ( .A(fanout_net_31 ), .B1(_02563_ ), .B2(_02564_ ), .ZN(_00877_ ) );
BUF_X8 _16244_ ( .A(_09471_ ), .Z(_02565_ ) );
BUF_X4 _16245_ ( .A(_02565_ ), .Z(_02566_ ) );
NAND4_X1 _16246_ ( .A1(_10267_ ), .A2(_02476_ ), .A3(_02472_ ), .A4(_02566_ ), .ZN(_02567_ ) );
OAI21_X1 _16247_ ( .A(\u_lsu.pmem[5925] ), .B1(_02474_ ), .B2(_02561_ ), .ZN(_02568_ ) );
AOI21_X1 _16248_ ( .A(fanout_net_31 ), .B1(_02567_ ), .B2(_02568_ ), .ZN(_00878_ ) );
AND2_X1 _16249_ ( .A1(_09141_ ), .A2(_02559_ ), .ZN(_02569_ ) );
OAI21_X1 _16250_ ( .A(_10715_ ), .B1(_02569_ ), .B2(\u_lsu.pmem[5924] ), .ZN(_02570_ ) );
AOI21_X1 _16251_ ( .A(_02570_ ), .B1(_09691_ ), .B2(_02569_ ), .ZN(_00879_ ) );
OAI21_X1 _16252_ ( .A(\u_lsu.pmem[5923] ), .B1(_02547_ ), .B2(_02561_ ), .ZN(_02571_ ) );
OR4_X1 _16253_ ( .A1(_09969_ ), .A2(_10042_ ), .A3(_02481_ ), .A4(_02560_ ), .ZN(_02572_ ) );
AOI21_X1 _16254_ ( .A(fanout_net_31 ), .B1(_02571_ ), .B2(_02572_ ), .ZN(_00880_ ) );
OAI21_X1 _16255_ ( .A(\u_lsu.pmem[5922] ), .B1(_02547_ ), .B2(_02561_ ), .ZN(_02573_ ) );
OR4_X1 _16256_ ( .A1(_09973_ ), .A2(_10042_ ), .A3(_02481_ ), .A4(_02560_ ), .ZN(_02574_ ) );
AOI21_X1 _16257_ ( .A(fanout_net_32 ), .B1(_02573_ ), .B2(_02574_ ), .ZN(_00881_ ) );
OAI21_X1 _16258_ ( .A(\u_lsu.pmem[5921] ), .B1(_02547_ ), .B2(_02561_ ), .ZN(_02575_ ) );
OR4_X1 _16259_ ( .A1(_09977_ ), .A2(_10042_ ), .A3(_02481_ ), .A4(_02560_ ), .ZN(_02576_ ) );
AOI21_X1 _16260_ ( .A(fanout_net_32 ), .B1(_02575_ ), .B2(_02576_ ), .ZN(_00882_ ) );
NAND4_X1 _16261_ ( .A1(_10279_ ), .A2(_02476_ ), .A3(_02472_ ), .A4(_02566_ ), .ZN(_02577_ ) );
OAI21_X1 _16262_ ( .A(\u_lsu.pmem[5920] ), .B1(_02474_ ), .B2(_02561_ ), .ZN(_02578_ ) );
AOI21_X1 _16263_ ( .A(fanout_net_32 ), .B1(_02577_ ), .B2(_02578_ ), .ZN(_00883_ ) );
NAND4_X1 _16264_ ( .A1(_10285_ ), .A2(_11039_ ), .A3(_02472_ ), .A4(_02566_ ), .ZN(_02579_ ) );
NAND3_X1 _16265_ ( .A1(_10289_ ), .A2(_02484_ ), .A3(_10286_ ), .ZN(_02580_ ) );
BUF_X4 _16266_ ( .A(_02580_ ), .Z(_02581_ ) );
OAI21_X1 _16267_ ( .A(\u_lsu.pmem[5895] ), .B1(_02474_ ), .B2(_02581_ ), .ZN(_02582_ ) );
AOI21_X1 _16268_ ( .A(fanout_net_32 ), .B1(_02579_ ), .B2(_02582_ ), .ZN(_00884_ ) );
NAND4_X1 _16269_ ( .A1(_10443_ ), .A2(_09713_ ), .A3(_02429_ ), .A4(_02371_ ), .ZN(_02583_ ) );
BUF_X4 _16270_ ( .A(_09730_ ), .Z(_02584_ ) );
OAI21_X1 _16271_ ( .A(\u_lsu.pmem[3717] ), .B1(_10425_ ), .B2(_02584_ ), .ZN(_02585_ ) );
AOI21_X1 _16272_ ( .A(fanout_net_32 ), .B1(_02583_ ), .B2(_02585_ ), .ZN(_00885_ ) );
NAND4_X1 _16273_ ( .A1(_10295_ ), .A2(_11039_ ), .A3(_02472_ ), .A4(_02566_ ), .ZN(_02586_ ) );
OAI21_X1 _16274_ ( .A(\u_lsu.pmem[5894] ), .B1(_02474_ ), .B2(_02581_ ), .ZN(_02587_ ) );
AOI21_X1 _16275_ ( .A(fanout_net_32 ), .B1(_02586_ ), .B2(_02587_ ), .ZN(_00886_ ) );
NAND4_X1 _16276_ ( .A1(_10299_ ), .A2(_11039_ ), .A3(_02472_ ), .A4(_02566_ ), .ZN(_02588_ ) );
OAI21_X1 _16277_ ( .A(\u_lsu.pmem[5893] ), .B1(_02474_ ), .B2(_02581_ ), .ZN(_02589_ ) );
AOI21_X1 _16278_ ( .A(fanout_net_32 ), .B1(_02588_ ), .B2(_02589_ ), .ZN(_00887_ ) );
NAND4_X1 _16279_ ( .A1(_10306_ ), .A2(_11039_ ), .A3(_02472_ ), .A4(_02566_ ), .ZN(_02590_ ) );
OAI21_X1 _16280_ ( .A(\u_lsu.pmem[5892] ), .B1(_02474_ ), .B2(_02581_ ), .ZN(_02591_ ) );
AOI21_X1 _16281_ ( .A(fanout_net_32 ), .B1(_02590_ ), .B2(_02591_ ), .ZN(_00888_ ) );
BUF_X4 _16282_ ( .A(_09673_ ), .Z(_02592_ ) );
NAND4_X1 _16283_ ( .A1(_10309_ ), .A2(_11039_ ), .A3(_02592_ ), .A4(_02566_ ), .ZN(_02593_ ) );
BUF_X4 _16284_ ( .A(_02209_ ), .Z(_02594_ ) );
OAI21_X1 _16285_ ( .A(\u_lsu.pmem[5891] ), .B1(_02594_ ), .B2(_02581_ ), .ZN(_02595_ ) );
AOI21_X1 _16286_ ( .A(fanout_net_32 ), .B1(_02593_ ), .B2(_02595_ ), .ZN(_00889_ ) );
OAI21_X1 _16287_ ( .A(\u_lsu.pmem[5890] ), .B1(_02547_ ), .B2(_02581_ ), .ZN(_02596_ ) );
NAND4_X1 _16288_ ( .A1(_09510_ ), .A2(_10976_ ), .A3(_09909_ ), .A4(_10313_ ), .ZN(_02597_ ) );
AOI21_X1 _16289_ ( .A(fanout_net_32 ), .B1(_02596_ ), .B2(_02597_ ), .ZN(_00890_ ) );
NAND4_X1 _16290_ ( .A1(_10316_ ), .A2(_11039_ ), .A3(_02592_ ), .A4(_02566_ ), .ZN(_02598_ ) );
OAI21_X1 _16291_ ( .A(\u_lsu.pmem[5889] ), .B1(_02594_ ), .B2(_02581_ ), .ZN(_02599_ ) );
AOI21_X1 _16292_ ( .A(fanout_net_32 ), .B1(_02598_ ), .B2(_02599_ ), .ZN(_00891_ ) );
BUF_X4 _16293_ ( .A(_10585_ ), .Z(_02600_ ) );
NAND4_X1 _16294_ ( .A1(_10320_ ), .A2(_02600_ ), .A3(_02592_ ), .A4(_02566_ ), .ZN(_02601_ ) );
OAI21_X1 _16295_ ( .A(\u_lsu.pmem[5888] ), .B1(_02594_ ), .B2(_02581_ ), .ZN(_02602_ ) );
AOI21_X1 _16296_ ( .A(fanout_net_32 ), .B1(_02601_ ), .B2(_02602_ ), .ZN(_00892_ ) );
NAND2_X1 _16297_ ( .A1(_09461_ ), .A2(_10324_ ), .ZN(_02603_ ) );
BUF_X4 _16298_ ( .A(_02603_ ), .Z(_02604_ ) );
OAI21_X1 _16299_ ( .A(\u_lsu.pmem[5863] ), .B1(_02547_ ), .B2(_02604_ ), .ZN(_02605_ ) );
NAND4_X1 _16300_ ( .A1(_02246_ ), .A2(_02382_ ), .A3(_09909_ ), .A4(_10324_ ), .ZN(_02606_ ) );
AOI21_X1 _16301_ ( .A(fanout_net_32 ), .B1(_02605_ ), .B2(_02606_ ), .ZN(_00893_ ) );
NAND4_X1 _16302_ ( .A1(_10332_ ), .A2(_02476_ ), .A3(_02592_ ), .A4(_02566_ ), .ZN(_02607_ ) );
OAI21_X1 _16303_ ( .A(\u_lsu.pmem[5862] ), .B1(_02594_ ), .B2(_02604_ ), .ZN(_02608_ ) );
AOI21_X1 _16304_ ( .A(fanout_net_32 ), .B1(_02607_ ), .B2(_02608_ ), .ZN(_00894_ ) );
BUF_X4 _16305_ ( .A(_02565_ ), .Z(_02609_ ) );
NAND4_X1 _16306_ ( .A1(_10336_ ), .A2(_02476_ ), .A3(_02592_ ), .A4(_02609_ ), .ZN(_02610_ ) );
OAI21_X1 _16307_ ( .A(\u_lsu.pmem[5861] ), .B1(_02594_ ), .B2(_02603_ ), .ZN(_02611_ ) );
AOI21_X1 _16308_ ( .A(fanout_net_32 ), .B1(_02610_ ), .B2(_02611_ ), .ZN(_00895_ ) );
NAND4_X1 _16309_ ( .A1(_10443_ ), .A2(_10453_ ), .A3(_02429_ ), .A4(_02371_ ), .ZN(_02612_ ) );
OAI21_X1 _16310_ ( .A(\u_lsu.pmem[3716] ), .B1(_10425_ ), .B2(_02584_ ), .ZN(_02613_ ) );
AOI21_X1 _16311_ ( .A(fanout_net_32 ), .B1(_02612_ ), .B2(_02613_ ), .ZN(_00896_ ) );
NAND4_X1 _16312_ ( .A1(_10339_ ), .A2(_02476_ ), .A3(_02592_ ), .A4(_02609_ ), .ZN(_02614_ ) );
OAI21_X1 _16313_ ( .A(\u_lsu.pmem[5860] ), .B1(_02594_ ), .B2(_02603_ ), .ZN(_02615_ ) );
AOI21_X1 _16314_ ( .A(fanout_net_32 ), .B1(_02614_ ), .B2(_02615_ ), .ZN(_00897_ ) );
NAND4_X1 _16315_ ( .A1(_10345_ ), .A2(_02476_ ), .A3(_02592_ ), .A4(_02609_ ), .ZN(_02616_ ) );
OAI21_X1 _16316_ ( .A(\u_lsu.pmem[5859] ), .B1(_02594_ ), .B2(_02603_ ), .ZN(_02617_ ) );
AOI21_X1 _16317_ ( .A(fanout_net_32 ), .B1(_02616_ ), .B2(_02617_ ), .ZN(_00898_ ) );
NAND4_X1 _16318_ ( .A1(_10350_ ), .A2(_02476_ ), .A3(_02592_ ), .A4(_02609_ ), .ZN(_02618_ ) );
OAI21_X1 _16319_ ( .A(\u_lsu.pmem[5858] ), .B1(_02594_ ), .B2(_02603_ ), .ZN(_02619_ ) );
AOI21_X1 _16320_ ( .A(fanout_net_32 ), .B1(_02618_ ), .B2(_02619_ ), .ZN(_00899_ ) );
BUF_X4 _16321_ ( .A(_10886_ ), .Z(_02620_ ) );
NAND4_X1 _16322_ ( .A1(_10354_ ), .A2(_02620_ ), .A3(_02592_ ), .A4(_02609_ ), .ZN(_02621_ ) );
OAI21_X1 _16323_ ( .A(\u_lsu.pmem[5857] ), .B1(_02594_ ), .B2(_02603_ ), .ZN(_02622_ ) );
AOI21_X1 _16324_ ( .A(fanout_net_32 ), .B1(_02621_ ), .B2(_02622_ ), .ZN(_00900_ ) );
NAND4_X1 _16325_ ( .A1(_10357_ ), .A2(_02620_ ), .A3(_02592_ ), .A4(_02609_ ), .ZN(_02623_ ) );
OAI21_X1 _16326_ ( .A(\u_lsu.pmem[5856] ), .B1(_02594_ ), .B2(_02603_ ), .ZN(_02624_ ) );
AOI21_X1 _16327_ ( .A(fanout_net_32 ), .B1(_02623_ ), .B2(_02624_ ), .ZN(_00901_ ) );
NAND2_X1 _16328_ ( .A1(_09461_ ), .A2(_10362_ ), .ZN(_02625_ ) );
BUF_X4 _16329_ ( .A(_02625_ ), .Z(_02626_ ) );
OAI21_X1 _16330_ ( .A(\u_lsu.pmem[5831] ), .B1(_02547_ ), .B2(_02626_ ), .ZN(_02627_ ) );
NAND4_X1 _16331_ ( .A1(_02246_ ), .A2(_02382_ ), .A3(_09909_ ), .A4(_10362_ ), .ZN(_02628_ ) );
AOI21_X1 _16332_ ( .A(fanout_net_32 ), .B1(_02627_ ), .B2(_02628_ ), .ZN(_00902_ ) );
BUF_X4 _16333_ ( .A(_09673_ ), .Z(_02629_ ) );
NAND4_X1 _16334_ ( .A1(_10368_ ), .A2(_02620_ ), .A3(_02629_ ), .A4(_02609_ ), .ZN(_02630_ ) );
BUF_X4 _16335_ ( .A(_02209_ ), .Z(_02631_ ) );
OAI21_X1 _16336_ ( .A(\u_lsu.pmem[5830] ), .B1(_02631_ ), .B2(_02626_ ), .ZN(_02632_ ) );
AOI21_X1 _16337_ ( .A(fanout_net_32 ), .B1(_02630_ ), .B2(_02632_ ), .ZN(_00903_ ) );
NAND4_X1 _16338_ ( .A1(_10371_ ), .A2(_02620_ ), .A3(_02629_ ), .A4(_02609_ ), .ZN(_02633_ ) );
OAI21_X1 _16339_ ( .A(\u_lsu.pmem[5829] ), .B1(_02631_ ), .B2(_02625_ ), .ZN(_02634_ ) );
AOI21_X1 _16340_ ( .A(fanout_net_32 ), .B1(_02633_ ), .B2(_02634_ ), .ZN(_00904_ ) );
NAND4_X1 _16341_ ( .A1(_10374_ ), .A2(_02620_ ), .A3(_02629_ ), .A4(_02609_ ), .ZN(_02635_ ) );
OAI21_X1 _16342_ ( .A(\u_lsu.pmem[5828] ), .B1(_02631_ ), .B2(_02625_ ), .ZN(_02636_ ) );
AOI21_X1 _16343_ ( .A(fanout_net_32 ), .B1(_02635_ ), .B2(_02636_ ), .ZN(_00905_ ) );
NAND4_X1 _16344_ ( .A1(_10377_ ), .A2(_02620_ ), .A3(_02629_ ), .A4(_02609_ ), .ZN(_02637_ ) );
OAI21_X1 _16345_ ( .A(\u_lsu.pmem[5827] ), .B1(_02631_ ), .B2(_02625_ ), .ZN(_02638_ ) );
AOI21_X1 _16346_ ( .A(fanout_net_32 ), .B1(_02637_ ), .B2(_02638_ ), .ZN(_00906_ ) );
NAND4_X1 _16347_ ( .A1(_10443_ ), .A2(_10456_ ), .A3(_02429_ ), .A4(_02371_ ), .ZN(_02639_ ) );
OAI21_X1 _16348_ ( .A(\u_lsu.pmem[3715] ), .B1(_10425_ ), .B2(_02584_ ), .ZN(_02640_ ) );
AOI21_X1 _16349_ ( .A(fanout_net_32 ), .B1(_02639_ ), .B2(_02640_ ), .ZN(_00907_ ) );
BUF_X4 _16350_ ( .A(_02565_ ), .Z(_02641_ ) );
NAND4_X1 _16351_ ( .A1(_10381_ ), .A2(_02620_ ), .A3(_02629_ ), .A4(_02641_ ), .ZN(_02642_ ) );
OAI21_X1 _16352_ ( .A(\u_lsu.pmem[5826] ), .B1(_02631_ ), .B2(_02625_ ), .ZN(_02643_ ) );
AOI21_X1 _16353_ ( .A(fanout_net_32 ), .B1(_02642_ ), .B2(_02643_ ), .ZN(_00908_ ) );
NAND4_X1 _16354_ ( .A1(_10384_ ), .A2(_02620_ ), .A3(_02629_ ), .A4(_02641_ ), .ZN(_02644_ ) );
OAI21_X1 _16355_ ( .A(\u_lsu.pmem[5825] ), .B1(_02631_ ), .B2(_02625_ ), .ZN(_02645_ ) );
AOI21_X1 _16356_ ( .A(fanout_net_32 ), .B1(_02644_ ), .B2(_02645_ ), .ZN(_00909_ ) );
NAND4_X1 _16357_ ( .A1(_10391_ ), .A2(_02620_ ), .A3(_02629_ ), .A4(_02641_ ), .ZN(_02646_ ) );
OAI21_X1 _16358_ ( .A(\u_lsu.pmem[5824] ), .B1(_02631_ ), .B2(_02625_ ), .ZN(_02647_ ) );
AOI21_X1 _16359_ ( .A(fanout_net_32 ), .B1(_02646_ ), .B2(_02647_ ), .ZN(_00910_ ) );
NAND4_X1 _16360_ ( .A1(_10394_ ), .A2(_02620_ ), .A3(_02629_ ), .A4(_02641_ ), .ZN(_02648_ ) );
NAND2_X1 _16361_ ( .A1(_09461_ ), .A2(_10398_ ), .ZN(_02649_ ) );
BUF_X4 _16362_ ( .A(_02649_ ), .Z(_02650_ ) );
OAI21_X1 _16363_ ( .A(\u_lsu.pmem[5799] ), .B1(_02631_ ), .B2(_02650_ ), .ZN(_02651_ ) );
AOI21_X1 _16364_ ( .A(fanout_net_33 ), .B1(_02648_ ), .B2(_02651_ ), .ZN(_00911_ ) );
BUF_X4 _16365_ ( .A(_10886_ ), .Z(_02652_ ) );
NAND4_X1 _16366_ ( .A1(_10402_ ), .A2(_02652_ ), .A3(_02629_ ), .A4(_02641_ ), .ZN(_02653_ ) );
OAI21_X1 _16367_ ( .A(\u_lsu.pmem[5798] ), .B1(_02631_ ), .B2(_02649_ ), .ZN(_02654_ ) );
AOI21_X1 _16368_ ( .A(fanout_net_33 ), .B1(_02653_ ), .B2(_02654_ ), .ZN(_00912_ ) );
NAND4_X1 _16369_ ( .A1(_10405_ ), .A2(_02652_ ), .A3(_02629_ ), .A4(_02641_ ), .ZN(_02655_ ) );
OAI21_X1 _16370_ ( .A(\u_lsu.pmem[5797] ), .B1(_02631_ ), .B2(_02649_ ), .ZN(_02656_ ) );
AOI21_X1 _16371_ ( .A(fanout_net_33 ), .B1(_02655_ ), .B2(_02656_ ), .ZN(_00913_ ) );
BUF_X8 _16372_ ( .A(_09455_ ), .Z(_02657_ ) );
BUF_X4 _16373_ ( .A(_02657_ ), .Z(_02658_ ) );
NAND4_X1 _16374_ ( .A1(_10408_ ), .A2(_02652_ ), .A3(_02658_ ), .A4(_02641_ ), .ZN(_02659_ ) );
BUF_X4 _16375_ ( .A(_02209_ ), .Z(_02660_ ) );
OAI21_X1 _16376_ ( .A(\u_lsu.pmem[5796] ), .B1(_02660_ ), .B2(_02649_ ), .ZN(_02661_ ) );
AOI21_X1 _16377_ ( .A(fanout_net_33 ), .B1(_02659_ ), .B2(_02661_ ), .ZN(_00914_ ) );
NAND4_X1 _16378_ ( .A1(_10411_ ), .A2(_02652_ ), .A3(_02658_ ), .A4(_02641_ ), .ZN(_02662_ ) );
OAI21_X1 _16379_ ( .A(\u_lsu.pmem[5795] ), .B1(_02660_ ), .B2(_02649_ ), .ZN(_02663_ ) );
AOI21_X1 _16380_ ( .A(fanout_net_33 ), .B1(_02662_ ), .B2(_02663_ ), .ZN(_00915_ ) );
NAND4_X1 _16381_ ( .A1(_10414_ ), .A2(_02652_ ), .A3(_02658_ ), .A4(_02641_ ), .ZN(_02664_ ) );
OAI21_X1 _16382_ ( .A(\u_lsu.pmem[5794] ), .B1(_02660_ ), .B2(_02649_ ), .ZN(_02665_ ) );
AOI21_X1 _16383_ ( .A(fanout_net_33 ), .B1(_02664_ ), .B2(_02665_ ), .ZN(_00916_ ) );
NAND4_X1 _16384_ ( .A1(_10417_ ), .A2(_02652_ ), .A3(_02658_ ), .A4(_02641_ ), .ZN(_02666_ ) );
OAI21_X1 _16385_ ( .A(\u_lsu.pmem[5793] ), .B1(_02660_ ), .B2(_02649_ ), .ZN(_02667_ ) );
AOI21_X1 _16386_ ( .A(fanout_net_33 ), .B1(_02666_ ), .B2(_02667_ ), .ZN(_00917_ ) );
BUF_X4 _16387_ ( .A(_02565_ ), .Z(_02668_ ) );
NAND4_X1 _16388_ ( .A1(_09775_ ), .A2(_02286_ ), .A3(_02658_ ), .A4(_02668_ ), .ZN(_02669_ ) );
OAI21_X1 _16389_ ( .A(\u_lsu.pmem[4323] ), .B1(_02660_ ), .B2(_09751_ ), .ZN(_02670_ ) );
AOI21_X1 _16390_ ( .A(fanout_net_33 ), .B1(_02669_ ), .B2(_02670_ ), .ZN(_00918_ ) );
OAI21_X1 _16391_ ( .A(\u_lsu.pmem[3714] ), .B1(_10426_ ), .B2(_09911_ ), .ZN(_02671_ ) );
BUF_X4 _16392_ ( .A(_11381_ ), .Z(_02672_ ) );
NAND4_X1 _16393_ ( .A1(_10460_ ), .A2(_10976_ ), .A3(_02672_ ), .A4(_02526_ ), .ZN(_02673_ ) );
AOI21_X1 _16394_ ( .A(fanout_net_33 ), .B1(_02671_ ), .B2(_02673_ ), .ZN(_00919_ ) );
BUF_X4 _16395_ ( .A(_11582_ ), .Z(_02674_ ) );
OAI21_X1 _16396_ ( .A(\u_lsu.pmem[5792] ), .B1(_02674_ ), .B2(_02650_ ), .ZN(_02675_ ) );
NAND4_X1 _16397_ ( .A1(_10525_ ), .A2(_02382_ ), .A3(_09909_ ), .A4(_10398_ ), .ZN(_02676_ ) );
AOI21_X1 _16398_ ( .A(fanout_net_33 ), .B1(_02675_ ), .B2(_02676_ ), .ZN(_00920_ ) );
NAND3_X1 _16399_ ( .A1(_10423_ ), .A2(_09875_ ), .A3(_09454_ ), .ZN(_02677_ ) );
BUF_X4 _16400_ ( .A(_02677_ ), .Z(_02678_ ) );
BUF_X4 _16401_ ( .A(_10901_ ), .Z(_02679_ ) );
OAI21_X1 _16402_ ( .A(\u_lsu.pmem[5767] ), .B1(_02678_ ), .B2(_02679_ ), .ZN(_02680_ ) );
NAND4_X1 _16403_ ( .A1(_10436_ ), .A2(_10976_ ), .A3(_09909_ ), .A4(_02345_ ), .ZN(_02681_ ) );
AOI21_X1 _16404_ ( .A(fanout_net_33 ), .B1(_02680_ ), .B2(_02681_ ), .ZN(_00921_ ) );
BUF_X4 _16405_ ( .A(_10442_ ), .Z(_02682_ ) );
NAND4_X1 _16406_ ( .A1(_02682_ ), .A2(_09658_ ), .A3(_02658_ ), .A4(_02668_ ), .ZN(_02683_ ) );
OAI21_X1 _16407_ ( .A(\u_lsu.pmem[5766] ), .B1(_02678_ ), .B2(_02492_ ), .ZN(_02684_ ) );
AOI21_X1 _16408_ ( .A(fanout_net_33 ), .B1(_02683_ ), .B2(_02684_ ), .ZN(_00922_ ) );
NAND4_X1 _16409_ ( .A1(_02682_ ), .A2(_09713_ ), .A3(_02658_ ), .A4(_02668_ ), .ZN(_02685_ ) );
OAI21_X1 _16410_ ( .A(\u_lsu.pmem[5765] ), .B1(_02678_ ), .B2(_02492_ ), .ZN(_02686_ ) );
AOI21_X1 _16411_ ( .A(fanout_net_33 ), .B1(_02685_ ), .B2(_02686_ ), .ZN(_00923_ ) );
NAND4_X1 _16412_ ( .A1(_02682_ ), .A2(_09514_ ), .A3(_02658_ ), .A4(_02668_ ), .ZN(_02687_ ) );
OAI21_X1 _16413_ ( .A(\u_lsu.pmem[5764] ), .B1(_02678_ ), .B2(_02492_ ), .ZN(_02688_ ) );
AOI21_X1 _16414_ ( .A(fanout_net_33 ), .B1(_02687_ ), .B2(_02688_ ), .ZN(_00924_ ) );
NAND4_X1 _16415_ ( .A1(_02682_ ), .A2(_10456_ ), .A3(_02658_ ), .A4(_02668_ ), .ZN(_02689_ ) );
OAI21_X1 _16416_ ( .A(\u_lsu.pmem[5763] ), .B1(_02678_ ), .B2(_02492_ ), .ZN(_02690_ ) );
AOI21_X1 _16417_ ( .A(fanout_net_33 ), .B1(_02689_ ), .B2(_02690_ ), .ZN(_00925_ ) );
OAI21_X1 _16418_ ( .A(\u_lsu.pmem[5762] ), .B1(_02678_ ), .B2(_02679_ ), .ZN(_02691_ ) );
NAND4_X1 _16419_ ( .A1(_10460_ ), .A2(_10976_ ), .A3(_09909_ ), .A4(_02345_ ), .ZN(_02692_ ) );
AOI21_X1 _16420_ ( .A(fanout_net_33 ), .B1(_02691_ ), .B2(_02692_ ), .ZN(_00926_ ) );
NAND4_X1 _16421_ ( .A1(_02682_ ), .A2(_09544_ ), .A3(_02658_ ), .A4(_02668_ ), .ZN(_02693_ ) );
BUF_X4 _16422_ ( .A(_09515_ ), .Z(_02694_ ) );
OAI21_X1 _16423_ ( .A(\u_lsu.pmem[5761] ), .B1(_02678_ ), .B2(_02694_ ), .ZN(_02695_ ) );
AOI21_X1 _16424_ ( .A(fanout_net_33 ), .B1(_02693_ ), .B2(_02695_ ), .ZN(_00927_ ) );
BUF_X4 _16425_ ( .A(_02657_ ), .Z(_02696_ ) );
NAND4_X1 _16426_ ( .A1(_02682_ ), .A2(_10467_ ), .A3(_02696_ ), .A4(_02668_ ), .ZN(_02697_ ) );
OAI21_X1 _16427_ ( .A(\u_lsu.pmem[5760] ), .B1(_02678_ ), .B2(_02694_ ), .ZN(_02698_ ) );
AOI21_X1 _16428_ ( .A(fanout_net_33 ), .B1(_02697_ ), .B2(_02698_ ), .ZN(_00928_ ) );
NAND2_X1 _16429_ ( .A1(_09475_ ), .A2(_10471_ ), .ZN(_02699_ ) );
BUF_X4 _16430_ ( .A(_02699_ ), .Z(_02700_ ) );
OAI21_X1 _16431_ ( .A(\u_lsu.pmem[5735] ), .B1(_02674_ ), .B2(_02700_ ), .ZN(_02701_ ) );
BUF_X4 _16432_ ( .A(_09476_ ), .Z(_02702_ ) );
NAND4_X1 _16433_ ( .A1(_02246_ ), .A2(_02382_ ), .A3(_02702_ ), .A4(_10489_ ), .ZN(_02703_ ) );
AOI21_X1 _16434_ ( .A(fanout_net_33 ), .B1(_02701_ ), .B2(_02703_ ), .ZN(_00929_ ) );
NAND4_X1 _16435_ ( .A1(_02682_ ), .A2(_09544_ ), .A3(_02429_ ), .A4(_02371_ ), .ZN(_02704_ ) );
OAI21_X1 _16436_ ( .A(\u_lsu.pmem[3713] ), .B1(_10425_ ), .B2(_02584_ ), .ZN(_02705_ ) );
AOI21_X1 _16437_ ( .A(fanout_net_33 ), .B1(_02704_ ), .B2(_02705_ ), .ZN(_00930_ ) );
OAI21_X1 _16438_ ( .A(\u_lsu.pmem[5734] ), .B1(_02674_ ), .B2(_02700_ ), .ZN(_02706_ ) );
NAND4_X1 _16439_ ( .A1(_11347_ ), .A2(_02382_ ), .A3(_02702_ ), .A4(_10489_ ), .ZN(_02707_ ) );
AOI21_X1 _16440_ ( .A(fanout_net_33 ), .B1(_02706_ ), .B2(_02707_ ), .ZN(_00931_ ) );
OAI21_X1 _16441_ ( .A(\u_lsu.pmem[5733] ), .B1(_02674_ ), .B2(_02699_ ), .ZN(_02708_ ) );
NAND4_X1 _16442_ ( .A1(_11351_ ), .A2(_02382_ ), .A3(_02702_ ), .A4(_10489_ ), .ZN(_02709_ ) );
AOI21_X1 _16443_ ( .A(fanout_net_33 ), .B1(_02708_ ), .B2(_02709_ ), .ZN(_00932_ ) );
OAI21_X1 _16444_ ( .A(\u_lsu.pmem[5732] ), .B1(_02674_ ), .B2(_02699_ ), .ZN(_02710_ ) );
NAND4_X1 _16445_ ( .A1(_02327_ ), .A2(_02382_ ), .A3(_02702_ ), .A4(_10489_ ), .ZN(_02711_ ) );
AOI21_X1 _16446_ ( .A(fanout_net_33 ), .B1(_02710_ ), .B2(_02711_ ), .ZN(_00933_ ) );
OAI21_X1 _16447_ ( .A(\u_lsu.pmem[5731] ), .B1(_02674_ ), .B2(_02699_ ), .ZN(_02712_ ) );
NAND4_X1 _16448_ ( .A1(_11385_ ), .A2(_02382_ ), .A3(_02702_ ), .A4(_10489_ ), .ZN(_02713_ ) );
AOI21_X1 _16449_ ( .A(fanout_net_33 ), .B1(_02712_ ), .B2(_02713_ ), .ZN(_00934_ ) );
OAI21_X1 _16450_ ( .A(\u_lsu.pmem[5730] ), .B1(_02674_ ), .B2(_02699_ ), .ZN(_02714_ ) );
NAND4_X1 _16451_ ( .A1(_02379_ ), .A2(_02382_ ), .A3(_02702_ ), .A4(_10489_ ), .ZN(_02715_ ) );
AOI21_X1 _16452_ ( .A(fanout_net_33 ), .B1(_02714_ ), .B2(_02715_ ), .ZN(_00935_ ) );
OAI21_X1 _16453_ ( .A(\u_lsu.pmem[5729] ), .B1(_02674_ ), .B2(_02699_ ), .ZN(_02716_ ) );
BUF_X4 _16454_ ( .A(_10548_ ), .Z(_02717_ ) );
NAND4_X1 _16455_ ( .A1(_11414_ ), .A2(_02717_ ), .A3(_02702_ ), .A4(_10471_ ), .ZN(_02718_ ) );
AOI21_X1 _16456_ ( .A(fanout_net_33 ), .B1(_02716_ ), .B2(_02718_ ), .ZN(_00936_ ) );
OAI21_X1 _16457_ ( .A(\u_lsu.pmem[5728] ), .B1(_02674_ ), .B2(_02699_ ), .ZN(_02719_ ) );
BUF_X4 _16458_ ( .A(_09621_ ), .Z(_02720_ ) );
NAND4_X1 _16459_ ( .A1(_02720_ ), .A2(_02717_ ), .A3(_02702_ ), .A4(_10471_ ), .ZN(_02721_ ) );
AOI21_X1 _16460_ ( .A(fanout_net_33 ), .B1(_02719_ ), .B2(_02721_ ), .ZN(_00937_ ) );
NAND2_X1 _16461_ ( .A1(_09475_ ), .A2(_10500_ ), .ZN(_02722_ ) );
BUF_X4 _16462_ ( .A(_02722_ ), .Z(_02723_ ) );
OAI21_X1 _16463_ ( .A(\u_lsu.pmem[5703] ), .B1(_02674_ ), .B2(_02723_ ), .ZN(_02724_ ) );
NAND4_X1 _16464_ ( .A1(_02246_ ), .A2(_02717_ ), .A3(_02702_ ), .A4(_10511_ ), .ZN(_02725_ ) );
AOI21_X1 _16465_ ( .A(fanout_net_33 ), .B1(_02724_ ), .B2(_02725_ ), .ZN(_00938_ ) );
BUF_X4 _16466_ ( .A(_11582_ ), .Z(_02726_ ) );
OAI21_X1 _16467_ ( .A(\u_lsu.pmem[5702] ), .B1(_02726_ ), .B2(_02723_ ), .ZN(_02727_ ) );
NAND4_X1 _16468_ ( .A1(_11347_ ), .A2(_02717_ ), .A3(_02702_ ), .A4(_10511_ ), .ZN(_02728_ ) );
AOI21_X1 _16469_ ( .A(fanout_net_33 ), .B1(_02727_ ), .B2(_02728_ ), .ZN(_00939_ ) );
OAI21_X1 _16470_ ( .A(\u_lsu.pmem[5701] ), .B1(_02726_ ), .B2(_02722_ ), .ZN(_02729_ ) );
BUF_X4 _16471_ ( .A(_09476_ ), .Z(_02730_ ) );
NAND4_X1 _16472_ ( .A1(_11351_ ), .A2(_02717_ ), .A3(_02730_ ), .A4(_10511_ ), .ZN(_02731_ ) );
AOI21_X1 _16473_ ( .A(fanout_net_33 ), .B1(_02729_ ), .B2(_02731_ ), .ZN(_00940_ ) );
NAND4_X1 _16474_ ( .A1(_02682_ ), .A2(_10467_ ), .A3(_02429_ ), .A4(_02371_ ), .ZN(_02732_ ) );
OAI21_X1 _16475_ ( .A(\u_lsu.pmem[3712] ), .B1(_10425_ ), .B2(_02584_ ), .ZN(_02733_ ) );
AOI21_X1 _16476_ ( .A(fanout_net_34 ), .B1(_02732_ ), .B2(_02733_ ), .ZN(_00941_ ) );
OAI21_X1 _16477_ ( .A(\u_lsu.pmem[5700] ), .B1(_02726_ ), .B2(_02722_ ), .ZN(_02734_ ) );
NAND4_X1 _16478_ ( .A1(_02327_ ), .A2(_02717_ ), .A3(_02730_ ), .A4(_10511_ ), .ZN(_02735_ ) );
AOI21_X1 _16479_ ( .A(fanout_net_34 ), .B1(_02734_ ), .B2(_02735_ ), .ZN(_00942_ ) );
OAI21_X1 _16480_ ( .A(\u_lsu.pmem[5699] ), .B1(_02726_ ), .B2(_02722_ ), .ZN(_02736_ ) );
NAND4_X1 _16481_ ( .A1(_11385_ ), .A2(_02717_ ), .A3(_02730_ ), .A4(_10500_ ), .ZN(_02737_ ) );
AOI21_X1 _16482_ ( .A(fanout_net_34 ), .B1(_02736_ ), .B2(_02737_ ), .ZN(_00943_ ) );
OAI21_X1 _16483_ ( .A(\u_lsu.pmem[5698] ), .B1(_02726_ ), .B2(_02722_ ), .ZN(_02738_ ) );
NAND4_X1 _16484_ ( .A1(_02379_ ), .A2(_02717_ ), .A3(_02730_ ), .A4(_10500_ ), .ZN(_02739_ ) );
AOI21_X1 _16485_ ( .A(fanout_net_34 ), .B1(_02738_ ), .B2(_02739_ ), .ZN(_00944_ ) );
OAI21_X1 _16486_ ( .A(\u_lsu.pmem[5697] ), .B1(_02726_ ), .B2(_02722_ ), .ZN(_02740_ ) );
NAND4_X1 _16487_ ( .A1(_11414_ ), .A2(_02717_ ), .A3(_02730_ ), .A4(_10500_ ), .ZN(_02741_ ) );
AOI21_X1 _16488_ ( .A(fanout_net_34 ), .B1(_02740_ ), .B2(_02741_ ), .ZN(_00945_ ) );
OAI21_X1 _16489_ ( .A(\u_lsu.pmem[5696] ), .B1(_02726_ ), .B2(_02722_ ), .ZN(_02742_ ) );
NAND4_X1 _16490_ ( .A1(_02720_ ), .A2(_02717_ ), .A3(_02730_ ), .A4(_10500_ ), .ZN(_02743_ ) );
AOI21_X1 _16491_ ( .A(fanout_net_34 ), .B1(_02742_ ), .B2(_02743_ ), .ZN(_00946_ ) );
NAND4_X1 _16492_ ( .A1(_10527_ ), .A2(_02652_ ), .A3(_02696_ ), .A4(_02668_ ), .ZN(_02744_ ) );
NAND2_X1 _16493_ ( .A1(_09475_ ), .A2(_10531_ ), .ZN(_02745_ ) );
OAI21_X1 _16494_ ( .A(\u_lsu.pmem[5671] ), .B1(_02660_ ), .B2(_02745_ ), .ZN(_02746_ ) );
AOI21_X1 _16495_ ( .A(fanout_net_34 ), .B1(_02744_ ), .B2(_02746_ ), .ZN(_00947_ ) );
NAND4_X1 _16496_ ( .A1(_10535_ ), .A2(_02652_ ), .A3(_02696_ ), .A4(_02668_ ), .ZN(_02747_ ) );
OAI21_X1 _16497_ ( .A(\u_lsu.pmem[5670] ), .B1(_02660_ ), .B2(_02745_ ), .ZN(_02748_ ) );
AOI21_X1 _16498_ ( .A(fanout_net_34 ), .B1(_02747_ ), .B2(_02748_ ), .ZN(_00948_ ) );
NAND4_X1 _16499_ ( .A1(_10538_ ), .A2(_02652_ ), .A3(_02696_ ), .A4(_02668_ ), .ZN(_02749_ ) );
OAI21_X1 _16500_ ( .A(\u_lsu.pmem[5669] ), .B1(_02660_ ), .B2(_02745_ ), .ZN(_02750_ ) );
AOI21_X1 _16501_ ( .A(fanout_net_34 ), .B1(_02749_ ), .B2(_02750_ ), .ZN(_00949_ ) );
BUF_X4 _16502_ ( .A(_02745_ ), .Z(_02751_ ) );
OAI21_X1 _16503_ ( .A(\u_lsu.pmem[5668] ), .B1(_02726_ ), .B2(_02751_ ), .ZN(_02752_ ) );
BUF_X4 _16504_ ( .A(_10548_ ), .Z(_02753_ ) );
NAND4_X1 _16505_ ( .A1(_02327_ ), .A2(_02753_ ), .A3(_02730_ ), .A4(_10542_ ), .ZN(_02754_ ) );
AOI21_X1 _16506_ ( .A(fanout_net_34 ), .B1(_02752_ ), .B2(_02754_ ), .ZN(_00950_ ) );
OAI21_X1 _16507_ ( .A(\u_lsu.pmem[5667] ), .B1(_02726_ ), .B2(_02751_ ), .ZN(_02755_ ) );
NAND4_X1 _16508_ ( .A1(_11385_ ), .A2(_02753_ ), .A3(_02730_ ), .A4(_10542_ ), .ZN(_02756_ ) );
AOI21_X1 _16509_ ( .A(fanout_net_34 ), .B1(_02755_ ), .B2(_02756_ ), .ZN(_00951_ ) );
BUF_X4 _16510_ ( .A(_10471_ ), .Z(_02757_ ) );
NAND4_X1 _16511_ ( .A1(_10018_ ), .A2(_11212_ ), .A3(_09914_ ), .A4(_02757_ ), .ZN(_02758_ ) );
OAI21_X1 _16512_ ( .A(\u_lsu.pmem[3687] ), .B1(_02342_ ), .B2(_10473_ ), .ZN(_02759_ ) );
AOI21_X1 _16513_ ( .A(fanout_net_34 ), .B1(_02758_ ), .B2(_02759_ ), .ZN(_00952_ ) );
OAI21_X1 _16514_ ( .A(\u_lsu.pmem[5666] ), .B1(_02726_ ), .B2(_02745_ ), .ZN(_02760_ ) );
NAND4_X1 _16515_ ( .A1(_02379_ ), .A2(_02753_ ), .A3(_02730_ ), .A4(_10531_ ), .ZN(_02761_ ) );
AOI21_X1 _16516_ ( .A(fanout_net_34 ), .B1(_02760_ ), .B2(_02761_ ), .ZN(_00953_ ) );
BUF_X4 _16517_ ( .A(_11582_ ), .Z(_02762_ ) );
OAI21_X1 _16518_ ( .A(\u_lsu.pmem[5665] ), .B1(_02762_ ), .B2(_02745_ ), .ZN(_02763_ ) );
NAND4_X1 _16519_ ( .A1(_11414_ ), .A2(_02753_ ), .A3(_02730_ ), .A4(_10531_ ), .ZN(_02764_ ) );
AOI21_X1 _16520_ ( .A(fanout_net_34 ), .B1(_02763_ ), .B2(_02764_ ), .ZN(_00954_ ) );
BUF_X4 _16521_ ( .A(_02565_ ), .Z(_02765_ ) );
NAND4_X1 _16522_ ( .A1(_10556_ ), .A2(_02652_ ), .A3(_02696_ ), .A4(_02765_ ), .ZN(_02766_ ) );
OAI21_X1 _16523_ ( .A(\u_lsu.pmem[5664] ), .B1(_02660_ ), .B2(_02745_ ), .ZN(_02767_ ) );
AOI21_X1 _16524_ ( .A(fanout_net_34 ), .B1(_02766_ ), .B2(_02767_ ), .ZN(_00955_ ) );
AND3_X1 _16525_ ( .A1(_10560_ ), .A2(_02409_ ), .A3(_10055_ ), .ZN(_02768_ ) );
INV_X1 _16526_ ( .A(_02768_ ), .ZN(_02769_ ) );
BUF_X4 _16527_ ( .A(_02769_ ), .Z(_02770_ ) );
OAI21_X1 _16528_ ( .A(\u_lsu.pmem[5639] ), .B1(_02762_ ), .B2(_02770_ ), .ZN(_02771_ ) );
BUF_X4 _16529_ ( .A(_02768_ ), .Z(_02772_ ) );
NAND3_X1 _16530_ ( .A1(_11139_ ), .A2(_11423_ ), .A3(_02772_ ), .ZN(_02773_ ) );
AOI21_X1 _16531_ ( .A(fanout_net_34 ), .B1(_02771_ ), .B2(_02773_ ), .ZN(_00956_ ) );
OAI21_X1 _16532_ ( .A(\u_lsu.pmem[5638] ), .B1(_02762_ ), .B2(_02770_ ), .ZN(_02774_ ) );
NAND3_X1 _16533_ ( .A1(_11139_ ), .A2(_10444_ ), .A3(_02772_ ), .ZN(_02775_ ) );
AOI21_X1 _16534_ ( .A(fanout_net_34 ), .B1(_02774_ ), .B2(_02775_ ), .ZN(_00957_ ) );
OAI21_X1 _16535_ ( .A(\u_lsu.pmem[5637] ), .B1(_02762_ ), .B2(_02770_ ), .ZN(_02776_ ) );
NAND3_X1 _16536_ ( .A1(_11139_ ), .A2(_10448_ ), .A3(_02772_ ), .ZN(_02777_ ) );
AOI21_X1 _16537_ ( .A(fanout_net_34 ), .B1(_02776_ ), .B2(_02777_ ), .ZN(_00958_ ) );
OAI21_X1 _16538_ ( .A(\u_lsu.pmem[5636] ), .B1(_02762_ ), .B2(_02770_ ), .ZN(_02778_ ) );
NAND3_X1 _16539_ ( .A1(_11139_ ), .A2(_10453_ ), .A3(_02772_ ), .ZN(_02779_ ) );
AOI21_X1 _16540_ ( .A(fanout_net_34 ), .B1(_02778_ ), .B2(_02779_ ), .ZN(_00959_ ) );
NAND4_X1 _16541_ ( .A1(_10575_ ), .A2(_02600_ ), .A3(_02696_ ), .A4(_02765_ ), .ZN(_02780_ ) );
OAI21_X1 _16542_ ( .A(\u_lsu.pmem[5635] ), .B1(_02660_ ), .B2(_02770_ ), .ZN(_02781_ ) );
AOI21_X1 _16543_ ( .A(fanout_net_34 ), .B1(_02780_ ), .B2(_02781_ ), .ZN(_00960_ ) );
NAND4_X1 _16544_ ( .A1(_10584_ ), .A2(_02486_ ), .A3(_10876_ ), .A4(_02765_ ), .ZN(_02782_ ) );
BUF_X4 _16545_ ( .A(_02209_ ), .Z(_02783_ ) );
OAI21_X1 _16546_ ( .A(\u_lsu.pmem[5634] ), .B1(_02783_ ), .B2(_02770_ ), .ZN(_02784_ ) );
AOI21_X1 _16547_ ( .A(fanout_net_34 ), .B1(_02782_ ), .B2(_02784_ ), .ZN(_00961_ ) );
OAI21_X1 _16548_ ( .A(\u_lsu.pmem[5633] ), .B1(_02762_ ), .B2(_02770_ ), .ZN(_02785_ ) );
NAND3_X1 _16549_ ( .A1(_11139_ ), .A2(_10463_ ), .A3(_02772_ ), .ZN(_02786_ ) );
AOI21_X1 _16550_ ( .A(fanout_net_34 ), .B1(_02785_ ), .B2(_02786_ ), .ZN(_00962_ ) );
NAND4_X1 _16551_ ( .A1(_10018_ ), .A2(_11212_ ), .A3(_09925_ ), .A4(_02757_ ), .ZN(_02787_ ) );
OAI21_X1 _16552_ ( .A(\u_lsu.pmem[3686] ), .B1(_02342_ ), .B2(_10473_ ), .ZN(_02788_ ) );
AOI21_X1 _16553_ ( .A(fanout_net_34 ), .B1(_02787_ ), .B2(_02788_ ), .ZN(_00963_ ) );
BUF_X4 _16554_ ( .A(_10886_ ), .Z(_02789_ ) );
NAND4_X1 _16555_ ( .A1(_10591_ ), .A2(_02789_ ), .A3(_02696_ ), .A4(_02765_ ), .ZN(_02790_ ) );
OAI21_X1 _16556_ ( .A(\u_lsu.pmem[5632] ), .B1(_02783_ ), .B2(_02770_ ), .ZN(_02791_ ) );
AOI21_X1 _16557_ ( .A(fanout_net_34 ), .B1(_02790_ ), .B2(_02791_ ), .ZN(_00964_ ) );
NAND2_X1 _16558_ ( .A1(_09461_ ), .A2(_10596_ ), .ZN(_02792_ ) );
BUF_X4 _16559_ ( .A(_02792_ ), .Z(_02793_ ) );
OAI21_X1 _16560_ ( .A(\u_lsu.pmem[5607] ), .B1(_02762_ ), .B2(_02793_ ), .ZN(_02794_ ) );
BUF_X4 _16561_ ( .A(_09476_ ), .Z(_02795_ ) );
NAND4_X1 _16562_ ( .A1(_02246_ ), .A2(_02753_ ), .A3(_02795_ ), .A4(_10596_ ), .ZN(_02796_ ) );
AOI21_X1 _16563_ ( .A(fanout_net_34 ), .B1(_02794_ ), .B2(_02796_ ), .ZN(_00965_ ) );
NAND4_X1 _16564_ ( .A1(_10603_ ), .A2(_02789_ ), .A3(_02696_ ), .A4(_02765_ ), .ZN(_02797_ ) );
OAI21_X1 _16565_ ( .A(\u_lsu.pmem[5606] ), .B1(_02783_ ), .B2(_02793_ ), .ZN(_02798_ ) );
AOI21_X1 _16566_ ( .A(fanout_net_34 ), .B1(_02797_ ), .B2(_02798_ ), .ZN(_00966_ ) );
NAND4_X1 _16567_ ( .A1(_10608_ ), .A2(_02600_ ), .A3(_02696_ ), .A4(_02765_ ), .ZN(_02799_ ) );
OAI21_X1 _16568_ ( .A(\u_lsu.pmem[5605] ), .B1(_02783_ ), .B2(_02792_ ), .ZN(_02800_ ) );
AOI21_X1 _16569_ ( .A(fanout_net_34 ), .B1(_02799_ ), .B2(_02800_ ), .ZN(_00967_ ) );
NAND4_X1 _16570_ ( .A1(_10611_ ), .A2(_02600_ ), .A3(_02696_ ), .A4(_02765_ ), .ZN(_02801_ ) );
OAI21_X1 _16571_ ( .A(\u_lsu.pmem[5604] ), .B1(_02783_ ), .B2(_02792_ ), .ZN(_02802_ ) );
AOI21_X1 _16572_ ( .A(fanout_net_34 ), .B1(_02801_ ), .B2(_02802_ ), .ZN(_00968_ ) );
BUF_X4 _16573_ ( .A(_02657_ ), .Z(_02803_ ) );
NAND4_X1 _16574_ ( .A1(_10614_ ), .A2(_02600_ ), .A3(_02803_ ), .A4(_02765_ ), .ZN(_02804_ ) );
OAI21_X1 _16575_ ( .A(\u_lsu.pmem[5603] ), .B1(_02783_ ), .B2(_02792_ ), .ZN(_02805_ ) );
AOI21_X1 _16576_ ( .A(fanout_net_34 ), .B1(_02804_ ), .B2(_02805_ ), .ZN(_00969_ ) );
NAND4_X1 _16577_ ( .A1(_10617_ ), .A2(_02600_ ), .A3(_02803_ ), .A4(_02765_ ), .ZN(_02806_ ) );
OAI21_X1 _16578_ ( .A(\u_lsu.pmem[5602] ), .B1(_02783_ ), .B2(_02792_ ), .ZN(_02807_ ) );
AOI21_X1 _16579_ ( .A(fanout_net_34 ), .B1(_02806_ ), .B2(_02807_ ), .ZN(_00970_ ) );
NAND4_X1 _16580_ ( .A1(_10621_ ), .A2(_02789_ ), .A3(_02803_ ), .A4(_02765_ ), .ZN(_02808_ ) );
OAI21_X1 _16581_ ( .A(\u_lsu.pmem[5601] ), .B1(_02783_ ), .B2(_02792_ ), .ZN(_02809_ ) );
AOI21_X1 _16582_ ( .A(fanout_net_35 ), .B1(_02808_ ), .B2(_02809_ ), .ZN(_00971_ ) );
BUF_X4 _16583_ ( .A(_02565_ ), .Z(_02810_ ) );
NAND4_X1 _16584_ ( .A1(_10624_ ), .A2(_02600_ ), .A3(_02803_ ), .A4(_02810_ ), .ZN(_02811_ ) );
OAI21_X1 _16585_ ( .A(\u_lsu.pmem[5600] ), .B1(_02783_ ), .B2(_02792_ ), .ZN(_02812_ ) );
AOI21_X1 _16586_ ( .A(fanout_net_35 ), .B1(_02811_ ), .B2(_02812_ ), .ZN(_00972_ ) );
NAND2_X1 _16587_ ( .A1(_09461_ ), .A2(_10627_ ), .ZN(_02813_ ) );
BUF_X4 _16588_ ( .A(_02813_ ), .Z(_02814_ ) );
OAI21_X1 _16589_ ( .A(\u_lsu.pmem[5575] ), .B1(_02762_ ), .B2(_02814_ ), .ZN(_02815_ ) );
NAND4_X1 _16590_ ( .A1(_02246_ ), .A2(_02753_ ), .A3(_02795_ ), .A4(_10627_ ), .ZN(_02816_ ) );
AOI21_X1 _16591_ ( .A(fanout_net_35 ), .B1(_02815_ ), .B2(_02816_ ), .ZN(_00973_ ) );
NAND4_X1 _16592_ ( .A1(_10018_ ), .A2(_11212_ ), .A3(_09928_ ), .A4(_02757_ ), .ZN(_02817_ ) );
OAI21_X1 _16593_ ( .A(\u_lsu.pmem[3685] ), .B1(_02342_ ), .B2(_10472_ ), .ZN(_02818_ ) );
AOI21_X1 _16594_ ( .A(fanout_net_35 ), .B1(_02817_ ), .B2(_02818_ ), .ZN(_00974_ ) );
NAND4_X1 _16595_ ( .A1(_10632_ ), .A2(_02600_ ), .A3(_02803_ ), .A4(_02810_ ), .ZN(_02819_ ) );
OAI21_X1 _16596_ ( .A(\u_lsu.pmem[5574] ), .B1(_02783_ ), .B2(_02814_ ), .ZN(_02820_ ) );
AOI21_X1 _16597_ ( .A(fanout_net_35 ), .B1(_02819_ ), .B2(_02820_ ), .ZN(_00975_ ) );
NAND4_X1 _16598_ ( .A1(_10635_ ), .A2(_02600_ ), .A3(_02803_ ), .A4(_02810_ ), .ZN(_02821_ ) );
BUF_X8 _16599_ ( .A(_09458_ ), .Z(_02822_ ) );
BUF_X4 _16600_ ( .A(_02822_ ), .Z(_02823_ ) );
OAI21_X1 _16601_ ( .A(\u_lsu.pmem[5573] ), .B1(_02823_ ), .B2(_02813_ ), .ZN(_02824_ ) );
AOI21_X1 _16602_ ( .A(fanout_net_35 ), .B1(_02821_ ), .B2(_02824_ ), .ZN(_00976_ ) );
NAND4_X1 _16603_ ( .A1(_10641_ ), .A2(_02600_ ), .A3(_02803_ ), .A4(_02810_ ), .ZN(_02825_ ) );
OAI21_X1 _16604_ ( .A(\u_lsu.pmem[5572] ), .B1(_02823_ ), .B2(_02813_ ), .ZN(_02826_ ) );
AOI21_X1 _16605_ ( .A(fanout_net_35 ), .B1(_02825_ ), .B2(_02826_ ), .ZN(_00977_ ) );
BUF_X4 _16606_ ( .A(_10585_ ), .Z(_02827_ ) );
NAND4_X1 _16607_ ( .A1(_10645_ ), .A2(_02827_ ), .A3(_02803_ ), .A4(_02810_ ), .ZN(_02828_ ) );
OAI21_X1 _16608_ ( .A(\u_lsu.pmem[5571] ), .B1(_02823_ ), .B2(_02813_ ), .ZN(_02829_ ) );
AOI21_X1 _16609_ ( .A(fanout_net_35 ), .B1(_02828_ ), .B2(_02829_ ), .ZN(_00978_ ) );
NAND4_X1 _16610_ ( .A1(_10649_ ), .A2(_02827_ ), .A3(_02803_ ), .A4(_02810_ ), .ZN(_02830_ ) );
OAI21_X1 _16611_ ( .A(\u_lsu.pmem[5570] ), .B1(_02823_ ), .B2(_02813_ ), .ZN(_02831_ ) );
AOI21_X1 _16612_ ( .A(fanout_net_35 ), .B1(_02830_ ), .B2(_02831_ ), .ZN(_00979_ ) );
NAND4_X1 _16613_ ( .A1(_10652_ ), .A2(_02789_ ), .A3(_02803_ ), .A4(_02810_ ), .ZN(_02832_ ) );
OAI21_X1 _16614_ ( .A(\u_lsu.pmem[5569] ), .B1(_02823_ ), .B2(_02813_ ), .ZN(_02833_ ) );
AOI21_X1 _16615_ ( .A(fanout_net_35 ), .B1(_02832_ ), .B2(_02833_ ), .ZN(_00980_ ) );
BUF_X4 _16616_ ( .A(_02657_ ), .Z(_02834_ ) );
NAND4_X1 _16617_ ( .A1(_10655_ ), .A2(_02827_ ), .A3(_02834_ ), .A4(_02810_ ), .ZN(_02835_ ) );
OAI21_X1 _16618_ ( .A(\u_lsu.pmem[5568] ), .B1(_02823_ ), .B2(_02813_ ), .ZN(_02836_ ) );
AOI21_X1 _16619_ ( .A(fanout_net_35 ), .B1(_02835_ ), .B2(_02836_ ), .ZN(_00981_ ) );
NAND4_X1 _16620_ ( .A1(_10658_ ), .A2(_02827_ ), .A3(_02834_ ), .A4(_02810_ ), .ZN(_02837_ ) );
NAND2_X1 _16621_ ( .A1(_09461_ ), .A2(_10661_ ), .ZN(_02838_ ) );
BUF_X4 _16622_ ( .A(_02838_ ), .Z(_02839_ ) );
OAI21_X1 _16623_ ( .A(\u_lsu.pmem[5543] ), .B1(_02823_ ), .B2(_02839_ ), .ZN(_02840_ ) );
AOI21_X1 _16624_ ( .A(fanout_net_35 ), .B1(_02837_ ), .B2(_02840_ ), .ZN(_00982_ ) );
NAND4_X1 _16625_ ( .A1(_10665_ ), .A2(_02789_ ), .A3(_02834_ ), .A4(_02810_ ), .ZN(_02841_ ) );
OAI21_X1 _16626_ ( .A(\u_lsu.pmem[5542] ), .B1(_02823_ ), .B2(_02838_ ), .ZN(_02842_ ) );
AOI21_X1 _16627_ ( .A(fanout_net_35 ), .B1(_02841_ ), .B2(_02842_ ), .ZN(_00983_ ) );
BUF_X4 _16628_ ( .A(_02565_ ), .Z(_02843_ ) );
NAND4_X1 _16629_ ( .A1(_10668_ ), .A2(_02827_ ), .A3(_02834_ ), .A4(_02843_ ), .ZN(_02844_ ) );
OAI21_X1 _16630_ ( .A(\u_lsu.pmem[5541] ), .B1(_02823_ ), .B2(_02838_ ), .ZN(_02845_ ) );
AOI21_X1 _16631_ ( .A(fanout_net_35 ), .B1(_02844_ ), .B2(_02845_ ), .ZN(_00984_ ) );
NAND4_X1 _16632_ ( .A1(_10018_ ), .A2(_11212_ ), .A3(_11151_ ), .A4(_02757_ ), .ZN(_02846_ ) );
OAI21_X1 _16633_ ( .A(\u_lsu.pmem[3684] ), .B1(_02342_ ), .B2(_10472_ ), .ZN(_02847_ ) );
AOI21_X1 _16634_ ( .A(fanout_net_35 ), .B1(_02846_ ), .B2(_02847_ ), .ZN(_00985_ ) );
NAND4_X1 _16635_ ( .A1(_10671_ ), .A2(_02789_ ), .A3(_02834_ ), .A4(_02843_ ), .ZN(_02848_ ) );
OAI21_X1 _16636_ ( .A(\u_lsu.pmem[5540] ), .B1(_02823_ ), .B2(_02838_ ), .ZN(_02849_ ) );
AOI21_X1 _16637_ ( .A(fanout_net_35 ), .B1(_02848_ ), .B2(_02849_ ), .ZN(_00986_ ) );
NAND4_X1 _16638_ ( .A1(_10674_ ), .A2(_02789_ ), .A3(_02834_ ), .A4(_02843_ ), .ZN(_02850_ ) );
BUF_X4 _16639_ ( .A(_02822_ ), .Z(_02851_ ) );
OAI21_X1 _16640_ ( .A(\u_lsu.pmem[5539] ), .B1(_02851_ ), .B2(_02838_ ), .ZN(_02852_ ) );
AOI21_X1 _16641_ ( .A(fanout_net_35 ), .B1(_02850_ ), .B2(_02852_ ), .ZN(_00987_ ) );
NAND4_X1 _16642_ ( .A1(_10679_ ), .A2(_02789_ ), .A3(_02834_ ), .A4(_02843_ ), .ZN(_02853_ ) );
OAI21_X1 _16643_ ( .A(\u_lsu.pmem[5538] ), .B1(_02851_ ), .B2(_02838_ ), .ZN(_02854_ ) );
AOI21_X1 _16644_ ( .A(fanout_net_35 ), .B1(_02853_ ), .B2(_02854_ ), .ZN(_00988_ ) );
NAND4_X1 _16645_ ( .A1(_10682_ ), .A2(_02789_ ), .A3(_02834_ ), .A4(_02843_ ), .ZN(_02855_ ) );
OAI21_X1 _16646_ ( .A(\u_lsu.pmem[5537] ), .B1(_02851_ ), .B2(_02838_ ), .ZN(_02856_ ) );
AOI21_X1 _16647_ ( .A(fanout_net_35 ), .B1(_02855_ ), .B2(_02856_ ), .ZN(_00989_ ) );
OAI21_X1 _16648_ ( .A(\u_lsu.pmem[5536] ), .B1(_02762_ ), .B2(_02839_ ), .ZN(_02857_ ) );
NAND4_X1 _16649_ ( .A1(_02720_ ), .A2(_02753_ ), .A3(_02795_ ), .A4(_10661_ ), .ZN(_02858_ ) );
AOI21_X1 _16650_ ( .A(fanout_net_35 ), .B1(_02857_ ), .B2(_02858_ ), .ZN(_00990_ ) );
NAND2_X1 _16651_ ( .A1(_10690_ ), .A2(_09475_ ), .ZN(_02859_ ) );
BUF_X4 _16652_ ( .A(_02859_ ), .Z(_02860_ ) );
OAI21_X1 _16653_ ( .A(\u_lsu.pmem[5511] ), .B1(_02860_ ), .B2(_02679_ ), .ZN(_02861_ ) );
BUF_X4 _16654_ ( .A(_10904_ ), .Z(_02862_ ) );
NAND4_X1 _16655_ ( .A1(_10695_ ), .A2(_10752_ ), .A3(_02795_ ), .A4(_02862_ ), .ZN(_02863_ ) );
AOI21_X1 _16656_ ( .A(fanout_net_35 ), .B1(_02861_ ), .B2(_02863_ ), .ZN(_00991_ ) );
OAI21_X1 _16657_ ( .A(\u_lsu.pmem[5510] ), .B1(_02860_ ), .B2(_02679_ ), .ZN(_02864_ ) );
NAND4_X1 _16658_ ( .A1(_10695_ ), .A2(_10185_ ), .A3(_02795_ ), .A4(_02862_ ), .ZN(_02865_ ) );
AOI21_X1 _16659_ ( .A(fanout_net_35 ), .B1(_02864_ ), .B2(_02865_ ), .ZN(_00992_ ) );
OAI21_X1 _16660_ ( .A(\u_lsu.pmem[5509] ), .B1(_02860_ ), .B2(_02679_ ), .ZN(_02866_ ) );
NAND4_X1 _16661_ ( .A1(_10695_ ), .A2(_10188_ ), .A3(_02795_ ), .A4(_02862_ ), .ZN(_02867_ ) );
AOI21_X1 _16662_ ( .A(fanout_net_35 ), .B1(_02866_ ), .B2(_02867_ ), .ZN(_00993_ ) );
OAI21_X1 _16663_ ( .A(\u_lsu.pmem[5508] ), .B1(_02860_ ), .B2(_02679_ ), .ZN(_02868_ ) );
BUF_X4 _16664_ ( .A(_10694_ ), .Z(_02869_ ) );
NAND4_X1 _16665_ ( .A1(_02869_ ), .A2(_10192_ ), .A3(_02795_ ), .A4(_02862_ ), .ZN(_02870_ ) );
AOI21_X1 _16666_ ( .A(fanout_net_35 ), .B1(_02868_ ), .B2(_02870_ ), .ZN(_00994_ ) );
OAI21_X1 _16667_ ( .A(\u_lsu.pmem[5507] ), .B1(_02860_ ), .B2(_02679_ ), .ZN(_02871_ ) );
NAND4_X1 _16668_ ( .A1(_02869_ ), .A2(_10915_ ), .A3(_02795_ ), .A4(_02862_ ), .ZN(_02872_ ) );
AOI21_X1 _16669_ ( .A(fanout_net_35 ), .B1(_02871_ ), .B2(_02872_ ), .ZN(_00995_ ) );
NAND4_X1 _16670_ ( .A1(_10018_ ), .A2(_11212_ ), .A3(_09934_ ), .A4(_02757_ ), .ZN(_02873_ ) );
BUF_X4 _16671_ ( .A(_09562_ ), .Z(_02874_ ) );
OAI21_X1 _16672_ ( .A(\u_lsu.pmem[3683] ), .B1(_02874_ ), .B2(_10472_ ), .ZN(_02875_ ) );
AOI21_X1 _16673_ ( .A(fanout_net_35 ), .B1(_02873_ ), .B2(_02875_ ), .ZN(_00996_ ) );
OAI21_X1 _16674_ ( .A(\u_lsu.pmem[5506] ), .B1(_02860_ ), .B2(_02679_ ), .ZN(_02876_ ) );
NAND4_X1 _16675_ ( .A1(_09537_ ), .A2(_10976_ ), .A3(_02795_ ), .A4(_02862_ ), .ZN(_02877_ ) );
AOI21_X1 _16676_ ( .A(fanout_net_35 ), .B1(_02876_ ), .B2(_02877_ ), .ZN(_00997_ ) );
OAI21_X1 _16677_ ( .A(\u_lsu.pmem[5505] ), .B1(_02860_ ), .B2(_02679_ ), .ZN(_02878_ ) );
NAND4_X1 _16678_ ( .A1(_02869_ ), .A2(_02308_ ), .A3(_02795_ ), .A4(_02862_ ), .ZN(_02879_ ) );
AOI21_X1 _16679_ ( .A(fanout_net_35 ), .B1(_02878_ ), .B2(_02879_ ), .ZN(_00998_ ) );
OAI21_X1 _16680_ ( .A(\u_lsu.pmem[5504] ), .B1(_02860_ ), .B2(_02679_ ), .ZN(_02880_ ) );
BUF_X8 _16681_ ( .A(_09475_ ), .Z(_02881_ ) );
BUF_X4 _16682_ ( .A(_02881_ ), .Z(_02882_ ) );
NAND4_X1 _16683_ ( .A1(_02869_ ), .A2(_11131_ ), .A3(_02882_ ), .A4(_02862_ ), .ZN(_02883_ ) );
AOI21_X1 _16684_ ( .A(fanout_net_35 ), .B1(_02880_ ), .B2(_02883_ ), .ZN(_00999_ ) );
AND3_X1 _16685_ ( .A1(_10055_ ), .A2(_02409_ ), .A3(_09558_ ), .ZN(_02884_ ) );
INV_X1 _16686_ ( .A(_02884_ ), .ZN(_02885_ ) );
NOR3_X1 _16687_ ( .A1(_09573_ ), .A2(_09741_ ), .A3(_02885_ ), .ZN(_02886_ ) );
AOI21_X1 _16688_ ( .A(\u_lsu.pmem[5479] ), .B1(_10182_ ), .B2(_02884_ ), .ZN(_02887_ ) );
NOR3_X1 _16689_ ( .A1(_02886_ ), .A2(fanout_net_35 ), .A3(_02887_ ), .ZN(_01000_ ) );
BUF_X4 _16690_ ( .A(_02885_ ), .Z(_02888_ ) );
OAI21_X1 _16691_ ( .A(\u_lsu.pmem[5478] ), .B1(_02762_ ), .B2(_02888_ ), .ZN(_02889_ ) );
NAND4_X1 _16692_ ( .A1(_11347_ ), .A2(_02753_ ), .A3(_02882_ ), .A4(_10723_ ), .ZN(_02890_ ) );
AOI21_X1 _16693_ ( .A(fanout_net_36 ), .B1(_02889_ ), .B2(_02890_ ), .ZN(_01001_ ) );
BUF_X4 _16694_ ( .A(_11582_ ), .Z(_02891_ ) );
OAI21_X1 _16695_ ( .A(\u_lsu.pmem[5477] ), .B1(_02891_ ), .B2(_02888_ ), .ZN(_02892_ ) );
NAND4_X1 _16696_ ( .A1(_11351_ ), .A2(_02753_ ), .A3(_02882_ ), .A4(_10723_ ), .ZN(_02893_ ) );
AOI21_X1 _16697_ ( .A(fanout_net_36 ), .B1(_02892_ ), .B2(_02893_ ), .ZN(_01002_ ) );
OAI21_X1 _16698_ ( .A(\u_lsu.pmem[5476] ), .B1(_02891_ ), .B2(_02888_ ), .ZN(_02894_ ) );
NAND4_X1 _16699_ ( .A1(_02327_ ), .A2(_02753_ ), .A3(_02882_ ), .A4(_10723_ ), .ZN(_02895_ ) );
AOI21_X1 _16700_ ( .A(fanout_net_36 ), .B1(_02894_ ), .B2(_02895_ ), .ZN(_01003_ ) );
OAI21_X1 _16701_ ( .A(\u_lsu.pmem[5475] ), .B1(_02891_ ), .B2(_02888_ ), .ZN(_02896_ ) );
BUF_X4 _16702_ ( .A(_10548_ ), .Z(_02897_ ) );
NAND4_X1 _16703_ ( .A1(_11385_ ), .A2(_02897_ ), .A3(_02882_ ), .A4(_10723_ ), .ZN(_02898_ ) );
AOI21_X1 _16704_ ( .A(fanout_net_36 ), .B1(_02896_ ), .B2(_02898_ ), .ZN(_01004_ ) );
OAI21_X1 _16705_ ( .A(\u_lsu.pmem[5474] ), .B1(_02891_ ), .B2(_02888_ ), .ZN(_02899_ ) );
NAND4_X1 _16706_ ( .A1(_02379_ ), .A2(_02897_ ), .A3(_02882_ ), .A4(_10723_ ), .ZN(_02900_ ) );
AOI21_X1 _16707_ ( .A(fanout_net_36 ), .B1(_02899_ ), .B2(_02900_ ), .ZN(_01005_ ) );
OAI21_X1 _16708_ ( .A(\u_lsu.pmem[5473] ), .B1(_02891_ ), .B2(_02888_ ), .ZN(_02901_ ) );
NAND4_X1 _16709_ ( .A1(_11414_ ), .A2(_02897_ ), .A3(_02882_ ), .A4(_10723_ ), .ZN(_02902_ ) );
AOI21_X1 _16710_ ( .A(fanout_net_36 ), .B1(_02901_ ), .B2(_02902_ ), .ZN(_01006_ ) );
BUF_X4 _16711_ ( .A(_09953_ ), .Z(_02903_ ) );
NAND4_X1 _16712_ ( .A1(_02903_ ), .A2(_11212_ ), .A3(_10015_ ), .A4(_02757_ ), .ZN(_02904_ ) );
OAI21_X1 _16713_ ( .A(\u_lsu.pmem[3682] ), .B1(_02874_ ), .B2(_10472_ ), .ZN(_02905_ ) );
AOI21_X1 _16714_ ( .A(fanout_net_36 ), .B1(_02904_ ), .B2(_02905_ ), .ZN(_01007_ ) );
OAI21_X1 _16715_ ( .A(\u_lsu.pmem[5472] ), .B1(_02891_ ), .B2(_02888_ ), .ZN(_02906_ ) );
NAND4_X1 _16716_ ( .A1(_02720_ ), .A2(_02897_ ), .A3(_02882_ ), .A4(_10723_ ), .ZN(_02907_ ) );
AOI21_X1 _16717_ ( .A(fanout_net_36 ), .B1(_02906_ ), .B2(_02907_ ), .ZN(_01008_ ) );
AND3_X1 _16718_ ( .A1(_10055_ ), .A2(_09020_ ), .A3(_09631_ ), .ZN(_02908_ ) );
INV_X1 _16719_ ( .A(_02908_ ), .ZN(_02909_ ) );
BUF_X4 _16720_ ( .A(_02909_ ), .Z(_02910_ ) );
OAI21_X1 _16721_ ( .A(\u_lsu.pmem[5447] ), .B1(_02891_ ), .B2(_02910_ ), .ZN(_02911_ ) );
OR4_X1 _16722_ ( .A1(_09565_ ), .A2(_10042_ ), .A3(_02481_ ), .A4(_02909_ ), .ZN(_02912_ ) );
AOI21_X1 _16723_ ( .A(fanout_net_36 ), .B1(_02911_ ), .B2(_02912_ ), .ZN(_01009_ ) );
OAI21_X1 _16724_ ( .A(\u_lsu.pmem[5446] ), .B1(_02891_ ), .B2(_02910_ ), .ZN(_02913_ ) );
NAND4_X1 _16725_ ( .A1(_11347_ ), .A2(_02897_ ), .A3(_02882_ ), .A4(_10750_ ), .ZN(_02914_ ) );
AOI21_X1 _16726_ ( .A(fanout_net_36 ), .B1(_02913_ ), .B2(_02914_ ), .ZN(_01010_ ) );
OAI21_X1 _16727_ ( .A(\u_lsu.pmem[5445] ), .B1(_02891_ ), .B2(_02910_ ), .ZN(_02915_ ) );
NAND4_X1 _16728_ ( .A1(_11351_ ), .A2(_02897_ ), .A3(_02882_ ), .A4(_10750_ ), .ZN(_02916_ ) );
AOI21_X1 _16729_ ( .A(fanout_net_36 ), .B1(_02915_ ), .B2(_02916_ ), .ZN(_01011_ ) );
OAI21_X1 _16730_ ( .A(\u_lsu.pmem[5444] ), .B1(_02891_ ), .B2(_02910_ ), .ZN(_02917_ ) );
BUF_X4 _16731_ ( .A(_02881_ ), .Z(_02918_ ) );
NAND4_X1 _16732_ ( .A1(_02327_ ), .A2(_02897_ ), .A3(_02918_ ), .A4(_10750_ ), .ZN(_02919_ ) );
AOI21_X1 _16733_ ( .A(fanout_net_36 ), .B1(_02917_ ), .B2(_02919_ ), .ZN(_01012_ ) );
BUF_X4 _16734_ ( .A(_11582_ ), .Z(_02920_ ) );
OAI21_X1 _16735_ ( .A(\u_lsu.pmem[5443] ), .B1(_02920_ ), .B2(_02910_ ), .ZN(_02921_ ) );
NAND4_X1 _16736_ ( .A1(_11385_ ), .A2(_02897_ ), .A3(_02918_ ), .A4(_10750_ ), .ZN(_02922_ ) );
AOI21_X1 _16737_ ( .A(fanout_net_36 ), .B1(_02921_ ), .B2(_02922_ ), .ZN(_01013_ ) );
OAI21_X1 _16738_ ( .A(\u_lsu.pmem[5442] ), .B1(_02920_ ), .B2(_02910_ ), .ZN(_02923_ ) );
NAND4_X1 _16739_ ( .A1(_02379_ ), .A2(_02897_ ), .A3(_02918_ ), .A4(_10750_ ), .ZN(_02924_ ) );
AOI21_X1 _16740_ ( .A(fanout_net_36 ), .B1(_02923_ ), .B2(_02924_ ), .ZN(_01014_ ) );
OAI21_X1 _16741_ ( .A(\u_lsu.pmem[5441] ), .B1(_02920_ ), .B2(_02910_ ), .ZN(_02925_ ) );
NAND4_X1 _16742_ ( .A1(_11414_ ), .A2(_02897_ ), .A3(_02918_ ), .A4(_10750_ ), .ZN(_02926_ ) );
AOI21_X1 _16743_ ( .A(fanout_net_36 ), .B1(_02925_ ), .B2(_02926_ ), .ZN(_01015_ ) );
OAI21_X1 _16744_ ( .A(\u_lsu.pmem[5440] ), .B1(_02920_ ), .B2(_02910_ ), .ZN(_02927_ ) );
BUF_X4 _16745_ ( .A(_09950_ ), .Z(_02928_ ) );
NAND4_X1 _16746_ ( .A1(_02720_ ), .A2(_02928_ ), .A3(_02918_ ), .A4(_10750_ ), .ZN(_02929_ ) );
AOI21_X1 _16747_ ( .A(fanout_net_36 ), .B1(_02927_ ), .B2(_02929_ ), .ZN(_01016_ ) );
NAND4_X1 _16748_ ( .A1(_09670_ ), .A2(_02789_ ), .A3(_02834_ ), .A4(_02843_ ), .ZN(_02930_ ) );
AND2_X2 _16749_ ( .A1(_09454_ ), .A2(_10773_ ), .ZN(_02931_ ) );
INV_X1 _16750_ ( .A(_02931_ ), .ZN(_02932_ ) );
BUF_X4 _16751_ ( .A(_02932_ ), .Z(_02933_ ) );
OAI21_X1 _16752_ ( .A(\u_lsu.pmem[5415] ), .B1(_02933_ ), .B2(_02694_ ), .ZN(_02934_ ) );
AOI21_X1 _16753_ ( .A(fanout_net_36 ), .B1(_02930_ ), .B2(_02934_ ), .ZN(_01017_ ) );
BUF_X4 _16754_ ( .A(_10065_ ), .Z(_02935_ ) );
NAND4_X1 _16755_ ( .A1(_02903_ ), .A2(_02935_ ), .A3(_09941_ ), .A4(_02757_ ), .ZN(_02936_ ) );
OAI21_X1 _16756_ ( .A(\u_lsu.pmem[3681] ), .B1(_02874_ ), .B2(_10472_ ), .ZN(_02937_ ) );
AOI21_X1 _16757_ ( .A(fanout_net_36 ), .B1(_02936_ ), .B2(_02937_ ), .ZN(_01018_ ) );
BUF_X4 _16758_ ( .A(_10886_ ), .Z(_02938_ ) );
NAND4_X1 _16759_ ( .A1(_09681_ ), .A2(_02938_ ), .A3(_02834_ ), .A4(_02843_ ), .ZN(_02939_ ) );
OAI21_X1 _16760_ ( .A(\u_lsu.pmem[5414] ), .B1(_02933_ ), .B2(_02694_ ), .ZN(_02940_ ) );
AOI21_X1 _16761_ ( .A(fanout_net_36 ), .B1(_02939_ ), .B2(_02940_ ), .ZN(_01019_ ) );
BUF_X4 _16762_ ( .A(_02657_ ), .Z(_02941_ ) );
NAND4_X1 _16763_ ( .A1(_09685_ ), .A2(_02938_ ), .A3(_02941_ ), .A4(_02843_ ), .ZN(_02942_ ) );
OAI21_X1 _16764_ ( .A(\u_lsu.pmem[5413] ), .B1(_02933_ ), .B2(_02694_ ), .ZN(_02943_ ) );
AOI21_X1 _16765_ ( .A(fanout_net_36 ), .B1(_02942_ ), .B2(_02943_ ), .ZN(_01020_ ) );
BUF_X4 _16766_ ( .A(_10901_ ), .Z(_02944_ ) );
OAI21_X1 _16767_ ( .A(\u_lsu.pmem[5412] ), .B1(_02933_ ), .B2(_02944_ ), .ZN(_02945_ ) );
NAND4_X1 _16768_ ( .A1(_02327_ ), .A2(_02928_ ), .A3(_02918_ ), .A4(_10773_ ), .ZN(_02946_ ) );
AOI21_X1 _16769_ ( .A(fanout_net_36 ), .B1(_02945_ ), .B2(_02946_ ), .ZN(_01021_ ) );
OAI21_X1 _16770_ ( .A(\u_lsu.pmem[5411] ), .B1(_02933_ ), .B2(_02944_ ), .ZN(_02947_ ) );
NAND4_X1 _16771_ ( .A1(_11385_ ), .A2(_02928_ ), .A3(_02918_ ), .A4(_10773_ ), .ZN(_02948_ ) );
AOI21_X1 _16772_ ( .A(fanout_net_36 ), .B1(_02947_ ), .B2(_02948_ ), .ZN(_01022_ ) );
OAI21_X1 _16773_ ( .A(\u_lsu.pmem[5410] ), .B1(_02933_ ), .B2(_02944_ ), .ZN(_02949_ ) );
NAND4_X1 _16774_ ( .A1(_02379_ ), .A2(_02928_ ), .A3(_02918_ ), .A4(_10773_ ), .ZN(_02950_ ) );
AOI21_X1 _16775_ ( .A(fanout_net_36 ), .B1(_02949_ ), .B2(_02950_ ), .ZN(_01023_ ) );
OAI21_X1 _16776_ ( .A(\u_lsu.pmem[5409] ), .B1(_02933_ ), .B2(_02944_ ), .ZN(_02951_ ) );
NAND4_X1 _16777_ ( .A1(_11414_ ), .A2(_02928_ ), .A3(_02918_ ), .A4(_10773_ ), .ZN(_02952_ ) );
AOI21_X1 _16778_ ( .A(fanout_net_36 ), .B1(_02951_ ), .B2(_02952_ ), .ZN(_01024_ ) );
NAND4_X1 _16779_ ( .A1(_09703_ ), .A2(_02938_ ), .A3(_02941_ ), .A4(_02843_ ), .ZN(_02953_ ) );
OAI21_X1 _16780_ ( .A(\u_lsu.pmem[5408] ), .B1(_02932_ ), .B2(_02694_ ), .ZN(_02954_ ) );
AOI21_X1 _16781_ ( .A(fanout_net_36 ), .B1(_02953_ ), .B2(_02954_ ), .ZN(_01025_ ) );
NAND4_X1 _16782_ ( .A1(_09708_ ), .A2(_02827_ ), .A3(_02941_ ), .A4(_02843_ ), .ZN(_02955_ ) );
NAND2_X1 _16783_ ( .A1(_09461_ ), .A2(_10797_ ), .ZN(_02956_ ) );
BUF_X4 _16784_ ( .A(_02956_ ), .Z(_02957_ ) );
OAI21_X1 _16785_ ( .A(\u_lsu.pmem[5383] ), .B1(_02851_ ), .B2(_02957_ ), .ZN(_02958_ ) );
AOI21_X1 _16786_ ( .A(fanout_net_36 ), .B1(_02955_ ), .B2(_02958_ ), .ZN(_01026_ ) );
BUF_X4 _16787_ ( .A(_02565_ ), .Z(_02959_ ) );
NAND4_X1 _16788_ ( .A1(_09715_ ), .A2(_02827_ ), .A3(_02941_ ), .A4(_02959_ ), .ZN(_02960_ ) );
OAI21_X1 _16789_ ( .A(\u_lsu.pmem[5382] ), .B1(_02851_ ), .B2(_02956_ ), .ZN(_02961_ ) );
AOI21_X1 _16790_ ( .A(fanout_net_36 ), .B1(_02960_ ), .B2(_02961_ ), .ZN(_01027_ ) );
NAND4_X1 _16791_ ( .A1(_09718_ ), .A2(_02827_ ), .A3(_02941_ ), .A4(_02959_ ), .ZN(_02962_ ) );
OAI21_X1 _16792_ ( .A(\u_lsu.pmem[5381] ), .B1(_02851_ ), .B2(_02956_ ), .ZN(_02963_ ) );
AOI21_X1 _16793_ ( .A(fanout_net_36 ), .B1(_02962_ ), .B2(_02963_ ), .ZN(_01028_ ) );
NAND4_X1 _16794_ ( .A1(_09780_ ), .A2(_02286_ ), .A3(_02941_ ), .A4(_02959_ ), .ZN(_02964_ ) );
OAI21_X1 _16795_ ( .A(\u_lsu.pmem[4322] ), .B1(_02851_ ), .B2(_09751_ ), .ZN(_02965_ ) );
AOI21_X1 _16796_ ( .A(fanout_net_36 ), .B1(_02964_ ), .B2(_02965_ ), .ZN(_01029_ ) );
NAND4_X1 _16797_ ( .A1(_02903_ ), .A2(_02935_ ), .A3(_09944_ ), .A4(_02757_ ), .ZN(_02966_ ) );
OAI21_X1 _16798_ ( .A(\u_lsu.pmem[3680] ), .B1(_02874_ ), .B2(_10472_ ), .ZN(_02967_ ) );
AOI21_X1 _16799_ ( .A(fanout_net_36 ), .B1(_02966_ ), .B2(_02967_ ), .ZN(_01030_ ) );
NAND4_X1 _16800_ ( .A1(_09721_ ), .A2(_02827_ ), .A3(_02941_ ), .A4(_02959_ ), .ZN(_02968_ ) );
OAI21_X1 _16801_ ( .A(\u_lsu.pmem[5380] ), .B1(_02851_ ), .B2(_02956_ ), .ZN(_02969_ ) );
AOI21_X1 _16802_ ( .A(fanout_net_37 ), .B1(_02968_ ), .B2(_02969_ ), .ZN(_01031_ ) );
NAND4_X1 _16803_ ( .A1(_09725_ ), .A2(_02827_ ), .A3(_02941_ ), .A4(_02959_ ), .ZN(_02970_ ) );
OAI21_X1 _16804_ ( .A(\u_lsu.pmem[5379] ), .B1(_02851_ ), .B2(_02956_ ), .ZN(_02971_ ) );
AOI21_X1 _16805_ ( .A(fanout_net_37 ), .B1(_02970_ ), .B2(_02971_ ), .ZN(_01032_ ) );
OAI21_X1 _16806_ ( .A(\u_lsu.pmem[5378] ), .B1(_02920_ ), .B2(_02957_ ), .ZN(_02972_ ) );
NAND4_X1 _16807_ ( .A1(_09510_ ), .A2(_09474_ ), .A3(_02918_ ), .A4(_10797_ ), .ZN(_02973_ ) );
AOI21_X1 _16808_ ( .A(fanout_net_37 ), .B1(_02972_ ), .B2(_02973_ ), .ZN(_01033_ ) );
NAND4_X1 _16809_ ( .A1(_09733_ ), .A2(_02938_ ), .A3(_02941_ ), .A4(_02959_ ), .ZN(_02974_ ) );
OAI21_X1 _16810_ ( .A(\u_lsu.pmem[5377] ), .B1(_02851_ ), .B2(_02956_ ), .ZN(_02975_ ) );
AOI21_X1 _16811_ ( .A(fanout_net_37 ), .B1(_02974_ ), .B2(_02975_ ), .ZN(_01034_ ) );
BUF_X4 _16812_ ( .A(_10585_ ), .Z(_02976_ ) );
NAND4_X1 _16813_ ( .A1(_09736_ ), .A2(_02976_ ), .A3(_02941_ ), .A4(_02959_ ), .ZN(_02977_ ) );
BUF_X4 _16814_ ( .A(_02822_ ), .Z(_02978_ ) );
OAI21_X1 _16815_ ( .A(\u_lsu.pmem[5376] ), .B1(_02978_ ), .B2(_02956_ ), .ZN(_02979_ ) );
AOI21_X1 _16816_ ( .A(fanout_net_37 ), .B1(_02977_ ), .B2(_02979_ ), .ZN(_01035_ ) );
BUF_X4 _16817_ ( .A(_09453_ ), .Z(_02980_ ) );
NAND2_X1 _16818_ ( .A1(_02980_ ), .A2(_10819_ ), .ZN(_02981_ ) );
BUF_X4 _16819_ ( .A(_02981_ ), .Z(_02982_ ) );
OAI21_X1 _16820_ ( .A(\u_lsu.pmem[5351] ), .B1(_02920_ ), .B2(_02982_ ), .ZN(_02983_ ) );
BUF_X4 _16821_ ( .A(_02881_ ), .Z(_02984_ ) );
NAND4_X1 _16822_ ( .A1(_02246_ ), .A2(_02928_ ), .A3(_02984_ ), .A4(_10819_ ), .ZN(_02985_ ) );
AOI21_X1 _16823_ ( .A(fanout_net_37 ), .B1(_02983_ ), .B2(_02985_ ), .ZN(_01036_ ) );
BUF_X4 _16824_ ( .A(_02657_ ), .Z(_02986_ ) );
NAND4_X1 _16825_ ( .A1(_09756_ ), .A2(_02976_ ), .A3(_02986_ ), .A4(_02959_ ), .ZN(_02987_ ) );
OAI21_X1 _16826_ ( .A(\u_lsu.pmem[5350] ), .B1(_02978_ ), .B2(_02982_ ), .ZN(_02988_ ) );
AOI21_X1 _16827_ ( .A(fanout_net_37 ), .B1(_02987_ ), .B2(_02988_ ), .ZN(_01037_ ) );
NAND4_X1 _16828_ ( .A1(_09763_ ), .A2(_02938_ ), .A3(_02986_ ), .A4(_02959_ ), .ZN(_02989_ ) );
OAI21_X1 _16829_ ( .A(\u_lsu.pmem[5349] ), .B1(_02978_ ), .B2(_02981_ ), .ZN(_02990_ ) );
AOI21_X1 _16830_ ( .A(fanout_net_37 ), .B1(_02989_ ), .B2(_02990_ ), .ZN(_01038_ ) );
NAND4_X1 _16831_ ( .A1(_09770_ ), .A2(_02976_ ), .A3(_02986_ ), .A4(_02959_ ), .ZN(_02991_ ) );
OAI21_X1 _16832_ ( .A(\u_lsu.pmem[5348] ), .B1(_02978_ ), .B2(_02981_ ), .ZN(_02992_ ) );
AOI21_X1 _16833_ ( .A(fanout_net_37 ), .B1(_02991_ ), .B2(_02992_ ), .ZN(_01039_ ) );
BUF_X4 _16834_ ( .A(_02565_ ), .Z(_02993_ ) );
NAND4_X1 _16835_ ( .A1(_09775_ ), .A2(_02938_ ), .A3(_02986_ ), .A4(_02993_ ), .ZN(_02994_ ) );
OAI21_X1 _16836_ ( .A(\u_lsu.pmem[5347] ), .B1(_02978_ ), .B2(_02981_ ), .ZN(_02995_ ) );
AOI21_X1 _16837_ ( .A(fanout_net_37 ), .B1(_02994_ ), .B2(_02995_ ), .ZN(_01040_ ) );
NOR2_X4 _16838_ ( .A1(_09450_ ), .A2(_10501_ ), .ZN(_02996_ ) );
NOR2_X1 _16839_ ( .A1(_02996_ ), .A2(\u_lsu.pmem[3655] ), .ZN(_02997_ ) );
AOI211_X1 _16840_ ( .A(fanout_net_37 ), .B(_02997_ ), .C1(_09568_ ), .C2(_02996_ ), .ZN(_01041_ ) );
NAND4_X1 _16841_ ( .A1(_09780_ ), .A2(_02938_ ), .A3(_02986_ ), .A4(_02993_ ), .ZN(_02998_ ) );
OAI21_X1 _16842_ ( .A(\u_lsu.pmem[5346] ), .B1(_02978_ ), .B2(_02981_ ), .ZN(_02999_ ) );
AOI21_X1 _16843_ ( .A(fanout_net_37 ), .B1(_02998_ ), .B2(_02999_ ), .ZN(_01042_ ) );
NAND4_X1 _16844_ ( .A1(_09787_ ), .A2(_02938_ ), .A3(_02986_ ), .A4(_02993_ ), .ZN(_03000_ ) );
OAI21_X1 _16845_ ( .A(\u_lsu.pmem[5345] ), .B1(_02978_ ), .B2(_02981_ ), .ZN(_03001_ ) );
AOI21_X1 _16846_ ( .A(fanout_net_37 ), .B1(_03000_ ), .B2(_03001_ ), .ZN(_01043_ ) );
NAND4_X1 _16847_ ( .A1(_09791_ ), .A2(_02938_ ), .A3(_02986_ ), .A4(_02993_ ), .ZN(_03002_ ) );
OAI21_X1 _16848_ ( .A(\u_lsu.pmem[5344] ), .B1(_02978_ ), .B2(_02981_ ), .ZN(_03003_ ) );
AOI21_X1 _16849_ ( .A(fanout_net_37 ), .B1(_03002_ ), .B2(_03003_ ), .ZN(_01044_ ) );
NAND2_X1 _16850_ ( .A1(_02980_ ), .A2(_10847_ ), .ZN(_03004_ ) );
BUF_X4 _16851_ ( .A(_03004_ ), .Z(_03005_ ) );
OAI21_X1 _16852_ ( .A(\u_lsu.pmem[5319] ), .B1(_02920_ ), .B2(_03005_ ), .ZN(_03006_ ) );
NAND4_X1 _16853_ ( .A1(_02246_ ), .A2(_02928_ ), .A3(_02984_ ), .A4(_10847_ ), .ZN(_03007_ ) );
AOI21_X1 _16854_ ( .A(fanout_net_37 ), .B1(_03006_ ), .B2(_03007_ ), .ZN(_01045_ ) );
NAND4_X1 _16855_ ( .A1(_09804_ ), .A2(_02486_ ), .A3(_10876_ ), .A4(_02993_ ), .ZN(_03008_ ) );
OAI21_X1 _16856_ ( .A(\u_lsu.pmem[5318] ), .B1(_02978_ ), .B2(_03005_ ), .ZN(_03009_ ) );
AOI21_X1 _16857_ ( .A(fanout_net_37 ), .B1(_03008_ ), .B2(_03009_ ), .ZN(_01046_ ) );
NAND4_X1 _16858_ ( .A1(_09811_ ), .A2(_02976_ ), .A3(_02986_ ), .A4(_02993_ ), .ZN(_03010_ ) );
OAI21_X1 _16859_ ( .A(\u_lsu.pmem[5317] ), .B1(_02978_ ), .B2(_03004_ ), .ZN(_03011_ ) );
AOI21_X1 _16860_ ( .A(fanout_net_37 ), .B1(_03010_ ), .B2(_03011_ ), .ZN(_01047_ ) );
NAND4_X1 _16861_ ( .A1(_09815_ ), .A2(_02976_ ), .A3(_02986_ ), .A4(_02993_ ), .ZN(_03012_ ) );
BUF_X4 _16862_ ( .A(_02822_ ), .Z(_03013_ ) );
OAI21_X1 _16863_ ( .A(\u_lsu.pmem[5316] ), .B1(_03013_ ), .B2(_03004_ ), .ZN(_03014_ ) );
AOI21_X1 _16864_ ( .A(fanout_net_37 ), .B1(_03012_ ), .B2(_03014_ ), .ZN(_01048_ ) );
NAND4_X1 _16865_ ( .A1(_09819_ ), .A2(_02976_ ), .A3(_02986_ ), .A4(_02993_ ), .ZN(_03015_ ) );
OAI21_X1 _16866_ ( .A(\u_lsu.pmem[5315] ), .B1(_03013_ ), .B2(_03004_ ), .ZN(_03016_ ) );
AOI21_X1 _16867_ ( .A(fanout_net_37 ), .B1(_03015_ ), .B2(_03016_ ), .ZN(_01049_ ) );
BUF_X4 _16868_ ( .A(_02657_ ), .Z(_03017_ ) );
NAND4_X1 _16869_ ( .A1(_09827_ ), .A2(_02938_ ), .A3(_03017_ ), .A4(_02993_ ), .ZN(_03018_ ) );
OAI21_X1 _16870_ ( .A(\u_lsu.pmem[5314] ), .B1(_03013_ ), .B2(_03004_ ), .ZN(_03019_ ) );
AOI21_X1 _16871_ ( .A(fanout_net_37 ), .B1(_03018_ ), .B2(_03019_ ), .ZN(_01050_ ) );
BUF_X8 _16872_ ( .A(_09875_ ), .Z(_03020_ ) );
BUF_X4 _16873_ ( .A(_03020_ ), .Z(_03021_ ) );
NAND4_X1 _16874_ ( .A1(_09831_ ), .A2(_03021_ ), .A3(_03017_ ), .A4(_02993_ ), .ZN(_03022_ ) );
OAI21_X1 _16875_ ( .A(\u_lsu.pmem[5313] ), .B1(_03013_ ), .B2(_03004_ ), .ZN(_03023_ ) );
AOI21_X1 _16876_ ( .A(fanout_net_37 ), .B1(_03022_ ), .B2(_03023_ ), .ZN(_01051_ ) );
NAND2_X1 _16877_ ( .A1(_02996_ ), .A2(_11145_ ), .ZN(_03024_ ) );
OAI21_X1 _16878_ ( .A(\u_lsu.pmem[3654] ), .B1(_02874_ ), .B2(_10502_ ), .ZN(_03025_ ) );
AOI21_X1 _16879_ ( .A(fanout_net_37 ), .B1(_03024_ ), .B2(_03025_ ), .ZN(_01052_ ) );
BUF_X4 _16880_ ( .A(_02565_ ), .Z(_03026_ ) );
NAND4_X1 _16881_ ( .A1(_09835_ ), .A2(_03021_ ), .A3(_03017_ ), .A4(_03026_ ), .ZN(_03027_ ) );
OAI21_X1 _16882_ ( .A(\u_lsu.pmem[5312] ), .B1(_03013_ ), .B2(_03004_ ), .ZN(_03028_ ) );
AOI21_X1 _16883_ ( .A(fanout_net_37 ), .B1(_03027_ ), .B2(_03028_ ), .ZN(_01053_ ) );
NAND4_X1 _16884_ ( .A1(_09840_ ), .A2(_03021_ ), .A3(_03017_ ), .A4(_03026_ ), .ZN(_03029_ ) );
NAND3_X1 _16885_ ( .A1(_09454_ ), .A2(_09743_ ), .A3(_09844_ ), .ZN(_03030_ ) );
BUF_X4 _16886_ ( .A(_03030_ ), .Z(_03031_ ) );
OAI21_X1 _16887_ ( .A(\u_lsu.pmem[5287] ), .B1(_03013_ ), .B2(_03031_ ), .ZN(_03032_ ) );
AOI21_X1 _16888_ ( .A(fanout_net_37 ), .B1(_03029_ ), .B2(_03032_ ), .ZN(_01054_ ) );
NAND4_X1 _16889_ ( .A1(_09849_ ), .A2(_02976_ ), .A3(_03017_ ), .A4(_03026_ ), .ZN(_03033_ ) );
OAI21_X1 _16890_ ( .A(\u_lsu.pmem[5286] ), .B1(_03013_ ), .B2(_03031_ ), .ZN(_03034_ ) );
AOI21_X1 _16891_ ( .A(fanout_net_37 ), .B1(_03033_ ), .B2(_03034_ ), .ZN(_01055_ ) );
NAND4_X1 _16892_ ( .A1(_09853_ ), .A2(_03021_ ), .A3(_03017_ ), .A4(_03026_ ), .ZN(_03035_ ) );
OAI21_X1 _16893_ ( .A(\u_lsu.pmem[5285] ), .B1(_03013_ ), .B2(_03030_ ), .ZN(_03036_ ) );
AOI21_X1 _16894_ ( .A(fanout_net_37 ), .B1(_03035_ ), .B2(_03036_ ), .ZN(_01056_ ) );
NAND4_X1 _16895_ ( .A1(_09858_ ), .A2(_03021_ ), .A3(_03017_ ), .A4(_03026_ ), .ZN(_03037_ ) );
OAI21_X1 _16896_ ( .A(\u_lsu.pmem[5284] ), .B1(_03013_ ), .B2(_03030_ ), .ZN(_03038_ ) );
AOI21_X1 _16897_ ( .A(fanout_net_37 ), .B1(_03037_ ), .B2(_03038_ ), .ZN(_01057_ ) );
NAND4_X1 _16898_ ( .A1(_09861_ ), .A2(_03021_ ), .A3(_03017_ ), .A4(_03026_ ), .ZN(_03039_ ) );
OAI21_X1 _16899_ ( .A(\u_lsu.pmem[5283] ), .B1(_03013_ ), .B2(_03030_ ), .ZN(_03040_ ) );
AOI21_X1 _16900_ ( .A(fanout_net_37 ), .B1(_03039_ ), .B2(_03040_ ), .ZN(_01058_ ) );
NAND4_X1 _16901_ ( .A1(_09864_ ), .A2(_03021_ ), .A3(_03017_ ), .A4(_03026_ ), .ZN(_03041_ ) );
BUF_X4 _16902_ ( .A(_02822_ ), .Z(_03042_ ) );
OAI21_X1 _16903_ ( .A(\u_lsu.pmem[5282] ), .B1(_03042_ ), .B2(_03030_ ), .ZN(_03043_ ) );
AOI21_X1 _16904_ ( .A(fanout_net_37 ), .B1(_03041_ ), .B2(_03043_ ), .ZN(_01059_ ) );
NAND4_X1 _16905_ ( .A1(_09867_ ), .A2(_03021_ ), .A3(_03017_ ), .A4(_03026_ ), .ZN(_03044_ ) );
OAI21_X1 _16906_ ( .A(\u_lsu.pmem[5281] ), .B1(_03042_ ), .B2(_03030_ ), .ZN(_03045_ ) );
AOI21_X1 _16907_ ( .A(fanout_net_37 ), .B1(_03044_ ), .B2(_03045_ ), .ZN(_01060_ ) );
BUF_X4 _16908_ ( .A(_02657_ ), .Z(_03046_ ) );
NAND4_X1 _16909_ ( .A1(_09881_ ), .A2(_02976_ ), .A3(_03046_ ), .A4(_03026_ ), .ZN(_03047_ ) );
OAI21_X1 _16910_ ( .A(\u_lsu.pmem[5280] ), .B1(_03042_ ), .B2(_03030_ ), .ZN(_03048_ ) );
AOI21_X1 _16911_ ( .A(fanout_net_38 ), .B1(_03047_ ), .B2(_03048_ ), .ZN(_01061_ ) );
OR3_X2 _16912_ ( .A1(_09889_ ), .A2(_09842_ ), .A3(_09135_ ), .ZN(_03049_ ) );
BUF_X4 _16913_ ( .A(_03049_ ), .Z(_03050_ ) );
OAI21_X1 _16914_ ( .A(\u_lsu.pmem[5255] ), .B1(_03050_ ), .B2(_02944_ ), .ZN(_03051_ ) );
NAND4_X1 _16915_ ( .A1(_10899_ ), .A2(_10752_ ), .A3(_02984_ ), .A4(_02862_ ), .ZN(_03052_ ) );
AOI21_X1 _16916_ ( .A(fanout_net_38 ), .B1(_03051_ ), .B2(_03052_ ), .ZN(_01062_ ) );
NAND2_X1 _16917_ ( .A1(_02996_ ), .A2(_11148_ ), .ZN(_03053_ ) );
OAI21_X1 _16918_ ( .A(\u_lsu.pmem[3653] ), .B1(_02874_ ), .B2(_10502_ ), .ZN(_03054_ ) );
AOI21_X1 _16919_ ( .A(fanout_net_38 ), .B1(_03053_ ), .B2(_03054_ ), .ZN(_01063_ ) );
OAI21_X1 _16920_ ( .A(\u_lsu.pmem[5254] ), .B1(_03050_ ), .B2(_02944_ ), .ZN(_03055_ ) );
BUF_X4 _16921_ ( .A(_09575_ ), .Z(_03056_ ) );
NAND4_X1 _16922_ ( .A1(_10899_ ), .A2(_03056_ ), .A3(_02984_ ), .A4(_02862_ ), .ZN(_03057_ ) );
AOI21_X1 _16923_ ( .A(fanout_net_38 ), .B1(_03055_ ), .B2(_03057_ ), .ZN(_01064_ ) );
OAI21_X1 _16924_ ( .A(\u_lsu.pmem[5253] ), .B1(_03050_ ), .B2(_02944_ ), .ZN(_03058_ ) );
BUF_X4 _16925_ ( .A(_09582_ ), .Z(_03059_ ) );
BUF_X4 _16926_ ( .A(_10904_ ), .Z(_03060_ ) );
NAND4_X1 _16927_ ( .A1(_10899_ ), .A2(_03059_ ), .A3(_02984_ ), .A4(_03060_ ), .ZN(_03061_ ) );
AOI21_X1 _16928_ ( .A(fanout_net_38 ), .B1(_03058_ ), .B2(_03061_ ), .ZN(_01065_ ) );
OAI21_X1 _16929_ ( .A(\u_lsu.pmem[5252] ), .B1(_03050_ ), .B2(_02944_ ), .ZN(_03062_ ) );
BUF_X4 _16930_ ( .A(_10898_ ), .Z(_03063_ ) );
BUF_X4 _16931_ ( .A(_08605_ ), .Z(_03064_ ) );
NAND4_X1 _16932_ ( .A1(_03063_ ), .A2(_03064_ ), .A3(_02984_ ), .A4(_03060_ ), .ZN(_03065_ ) );
AOI21_X1 _16933_ ( .A(fanout_net_38 ), .B1(_03062_ ), .B2(_03065_ ), .ZN(_01066_ ) );
OAI21_X1 _16934_ ( .A(\u_lsu.pmem[5251] ), .B1(_03050_ ), .B2(_02944_ ), .ZN(_03066_ ) );
NAND4_X1 _16935_ ( .A1(_03063_ ), .A2(_10915_ ), .A3(_02984_ ), .A4(_03060_ ), .ZN(_03067_ ) );
AOI21_X1 _16936_ ( .A(fanout_net_38 ), .B1(_03066_ ), .B2(_03067_ ), .ZN(_01067_ ) );
OAI21_X1 _16937_ ( .A(\u_lsu.pmem[5250] ), .B1(_03050_ ), .B2(_02944_ ), .ZN(_03068_ ) );
NAND4_X1 _16938_ ( .A1(_09906_ ), .A2(_10976_ ), .A3(_02984_ ), .A4(_03060_ ), .ZN(_03069_ ) );
AOI21_X1 _16939_ ( .A(fanout_net_38 ), .B1(_03068_ ), .B2(_03069_ ), .ZN(_01068_ ) );
BUF_X4 _16940_ ( .A(_10901_ ), .Z(_03070_ ) );
OAI21_X1 _16941_ ( .A(\u_lsu.pmem[5249] ), .B1(_03050_ ), .B2(_03070_ ), .ZN(_03071_ ) );
NAND4_X1 _16942_ ( .A1(_03063_ ), .A2(_02308_ ), .A3(_02984_ ), .A4(_03060_ ), .ZN(_03072_ ) );
AOI21_X1 _16943_ ( .A(fanout_net_38 ), .B1(_03071_ ), .B2(_03072_ ), .ZN(_01069_ ) );
OAI21_X1 _16944_ ( .A(\u_lsu.pmem[5248] ), .B1(_03050_ ), .B2(_03070_ ), .ZN(_03073_ ) );
NAND4_X1 _16945_ ( .A1(_03063_ ), .A2(_11131_ ), .A3(_02984_ ), .A4(_03060_ ), .ZN(_03074_ ) );
AOI21_X1 _16946_ ( .A(fanout_net_38 ), .B1(_03073_ ), .B2(_03074_ ), .ZN(_01070_ ) );
NAND3_X1 _16947_ ( .A1(_09915_ ), .A2(_09743_ ), .A3(_02409_ ), .ZN(_03075_ ) );
BUF_X4 _16948_ ( .A(_03075_ ), .Z(_03076_ ) );
OAI21_X1 _16949_ ( .A(\u_lsu.pmem[5223] ), .B1(_02920_ ), .B2(_03076_ ), .ZN(_03077_ ) );
OR4_X1 _16950_ ( .A1(_09565_ ), .A2(_03075_ ), .A3(_02481_ ), .A4(_09498_ ), .ZN(_03078_ ) );
AOI21_X1 _16951_ ( .A(fanout_net_38 ), .B1(_03077_ ), .B2(_03078_ ), .ZN(_01071_ ) );
OAI21_X1 _16952_ ( .A(\u_lsu.pmem[5222] ), .B1(_02920_ ), .B2(_03076_ ), .ZN(_03079_ ) );
BUF_X4 _16953_ ( .A(_02881_ ), .Z(_03080_ ) );
NAND4_X1 _16954_ ( .A1(_11347_ ), .A2(_02928_ ), .A3(_03080_ ), .A4(_10939_ ), .ZN(_03081_ ) );
AOI21_X1 _16955_ ( .A(fanout_net_38 ), .B1(_03079_ ), .B2(_03081_ ), .ZN(_01072_ ) );
OAI21_X1 _16956_ ( .A(\u_lsu.pmem[5221] ), .B1(_02920_ ), .B2(_03076_ ), .ZN(_03082_ ) );
NAND4_X1 _16957_ ( .A1(_11351_ ), .A2(_02928_ ), .A3(_03080_ ), .A4(_10939_ ), .ZN(_03083_ ) );
AOI21_X1 _16958_ ( .A(fanout_net_38 ), .B1(_03082_ ), .B2(_03083_ ), .ZN(_01073_ ) );
BUF_X4 _16959_ ( .A(_11151_ ), .Z(_03084_ ) );
NAND2_X1 _16960_ ( .A1(_02996_ ), .A2(_03084_ ), .ZN(_03085_ ) );
OAI21_X1 _16961_ ( .A(\u_lsu.pmem[3652] ), .B1(_02874_ ), .B2(_10501_ ), .ZN(_03086_ ) );
AOI21_X1 _16962_ ( .A(fanout_net_38 ), .B1(_03085_ ), .B2(_03086_ ), .ZN(_01074_ ) );
BUF_X4 _16963_ ( .A(_09459_ ), .Z(_03087_ ) );
OAI21_X1 _16964_ ( .A(\u_lsu.pmem[5220] ), .B1(_03087_ ), .B2(_03076_ ), .ZN(_03088_ ) );
NAND4_X1 _16965_ ( .A1(_02327_ ), .A2(_02928_ ), .A3(_03080_ ), .A4(_10939_ ), .ZN(_03089_ ) );
AOI21_X1 _16966_ ( .A(fanout_net_38 ), .B1(_03088_ ), .B2(_03089_ ), .ZN(_01075_ ) );
OAI21_X1 _16967_ ( .A(\u_lsu.pmem[5219] ), .B1(_03087_ ), .B2(_03076_ ), .ZN(_03090_ ) );
BUF_X4 _16968_ ( .A(_09448_ ), .Z(_03091_ ) );
BUF_X4 _16969_ ( .A(_09950_ ), .Z(_03092_ ) );
NAND4_X1 _16970_ ( .A1(_03091_ ), .A2(_03092_ ), .A3(_03080_ ), .A4(_10939_ ), .ZN(_03093_ ) );
AOI21_X1 _16971_ ( .A(fanout_net_38 ), .B1(_03090_ ), .B2(_03093_ ), .ZN(_01076_ ) );
OAI21_X1 _16972_ ( .A(\u_lsu.pmem[5218] ), .B1(_03087_ ), .B2(_03076_ ), .ZN(_03094_ ) );
NAND4_X1 _16973_ ( .A1(_02379_ ), .A2(_03092_ ), .A3(_03080_ ), .A4(_10939_ ), .ZN(_03095_ ) );
AOI21_X1 _16974_ ( .A(fanout_net_38 ), .B1(_03094_ ), .B2(_03095_ ), .ZN(_01077_ ) );
OAI21_X1 _16975_ ( .A(\u_lsu.pmem[5217] ), .B1(_03087_ ), .B2(_03076_ ), .ZN(_03096_ ) );
NAND4_X1 _16976_ ( .A1(_11414_ ), .A2(_03092_ ), .A3(_03080_ ), .A4(_10929_ ), .ZN(_03097_ ) );
AOI21_X1 _16977_ ( .A(fanout_net_38 ), .B1(_03096_ ), .B2(_03097_ ), .ZN(_01078_ ) );
OAI21_X1 _16978_ ( .A(\u_lsu.pmem[5216] ), .B1(_03087_ ), .B2(_03076_ ), .ZN(_03098_ ) );
NAND4_X1 _16979_ ( .A1(_02720_ ), .A2(_03092_ ), .A3(_03080_ ), .A4(_10929_ ), .ZN(_03099_ ) );
AOI21_X1 _16980_ ( .A(fanout_net_38 ), .B1(_03098_ ), .B2(_03099_ ), .ZN(_01079_ ) );
NAND3_X1 _16981_ ( .A1(_09948_ ), .A2(_02409_ ), .A3(_10286_ ), .ZN(_03100_ ) );
BUF_X4 _16982_ ( .A(_03100_ ), .Z(_03101_ ) );
OAI21_X1 _16983_ ( .A(\u_lsu.pmem[5191] ), .B1(_03087_ ), .B2(_03101_ ), .ZN(_03102_ ) );
OR4_X1 _16984_ ( .A1(_09565_ ), .A2(_03100_ ), .A3(_02481_ ), .A4(_09498_ ), .ZN(_03103_ ) );
AOI21_X1 _16985_ ( .A(fanout_net_38 ), .B1(_03102_ ), .B2(_03103_ ), .ZN(_01080_ ) );
OAI21_X1 _16986_ ( .A(\u_lsu.pmem[5190] ), .B1(_03087_ ), .B2(_03101_ ), .ZN(_03104_ ) );
NAND4_X1 _16987_ ( .A1(_09957_ ), .A2(_10976_ ), .A3(_03080_ ), .A4(_03060_ ), .ZN(_03105_ ) );
AOI21_X1 _16988_ ( .A(fanout_net_38 ), .B1(_03104_ ), .B2(_03105_ ), .ZN(_01081_ ) );
OAI21_X1 _16989_ ( .A(\u_lsu.pmem[5189] ), .B1(_03087_ ), .B2(_03101_ ), .ZN(_03106_ ) );
BUF_X4 _16990_ ( .A(_10063_ ), .Z(_03107_ ) );
NAND4_X1 _16991_ ( .A1(_09961_ ), .A2(_03107_ ), .A3(_03080_ ), .A4(_03060_ ), .ZN(_03108_ ) );
AOI21_X1 _16992_ ( .A(fanout_net_38 ), .B1(_03106_ ), .B2(_03108_ ), .ZN(_01082_ ) );
OAI21_X1 _16993_ ( .A(\u_lsu.pmem[5188] ), .B1(_03087_ ), .B2(_03101_ ), .ZN(_03109_ ) );
NAND4_X1 _16994_ ( .A1(_09966_ ), .A2(_03107_ ), .A3(_03080_ ), .A4(_03060_ ), .ZN(_03110_ ) );
AOI21_X1 _16995_ ( .A(fanout_net_38 ), .B1(_03109_ ), .B2(_03110_ ), .ZN(_01083_ ) );
OAI21_X1 _16996_ ( .A(\u_lsu.pmem[5187] ), .B1(_03087_ ), .B2(_03101_ ), .ZN(_03111_ ) );
BUF_X4 _16997_ ( .A(_02881_ ), .Z(_03112_ ) );
NAND4_X1 _16998_ ( .A1(_09970_ ), .A2(_03107_ ), .A3(_03112_ ), .A4(_03060_ ), .ZN(_03113_ ) );
AOI21_X1 _16999_ ( .A(fanout_net_38 ), .B1(_03111_ ), .B2(_03113_ ), .ZN(_01084_ ) );
BUF_X4 _17000_ ( .A(_09448_ ), .Z(_03114_ ) );
NAND2_X1 _17001_ ( .A1(_02996_ ), .A2(_03114_ ), .ZN(_03115_ ) );
OAI21_X1 _17002_ ( .A(\u_lsu.pmem[3651] ), .B1(_02874_ ), .B2(_10501_ ), .ZN(_03116_ ) );
AOI21_X1 _17003_ ( .A(fanout_net_38 ), .B1(_03115_ ), .B2(_03116_ ), .ZN(_01085_ ) );
BUF_X4 _17004_ ( .A(_09459_ ), .Z(_03117_ ) );
OAI21_X1 _17005_ ( .A(\u_lsu.pmem[5186] ), .B1(_03117_ ), .B2(_03101_ ), .ZN(_03118_ ) );
BUF_X4 _17006_ ( .A(_10904_ ), .Z(_03119_ ) );
NAND4_X1 _17007_ ( .A1(_09974_ ), .A2(_03107_ ), .A3(_03112_ ), .A4(_03119_ ), .ZN(_03120_ ) );
AOI21_X1 _17008_ ( .A(fanout_net_38 ), .B1(_03118_ ), .B2(_03120_ ), .ZN(_01086_ ) );
OAI21_X1 _17009_ ( .A(\u_lsu.pmem[5185] ), .B1(_03117_ ), .B2(_03101_ ), .ZN(_03121_ ) );
NAND4_X1 _17010_ ( .A1(_09978_ ), .A2(_03107_ ), .A3(_03112_ ), .A4(_03119_ ), .ZN(_03122_ ) );
AOI21_X1 _17011_ ( .A(fanout_net_38 ), .B1(_03121_ ), .B2(_03122_ ), .ZN(_01087_ ) );
OAI21_X1 _17012_ ( .A(\u_lsu.pmem[5184] ), .B1(_03117_ ), .B2(_03101_ ), .ZN(_03123_ ) );
NAND4_X1 _17013_ ( .A1(_09982_ ), .A2(_03107_ ), .A3(_03112_ ), .A4(_03119_ ), .ZN(_03124_ ) );
AOI21_X1 _17014_ ( .A(fanout_net_38 ), .B1(_03123_ ), .B2(_03124_ ), .ZN(_01088_ ) );
NAND4_X1 _17015_ ( .A1(_09987_ ), .A2(_03021_ ), .A3(_03046_ ), .A4(_03026_ ), .ZN(_03125_ ) );
NAND3_X1 _17016_ ( .A1(_09989_ ), .A2(_09743_ ), .A3(_02484_ ), .ZN(_03126_ ) );
BUF_X4 _17017_ ( .A(_03126_ ), .Z(_03127_ ) );
OAI21_X1 _17018_ ( .A(\u_lsu.pmem[5159] ), .B1(_03042_ ), .B2(_03127_ ), .ZN(_03128_ ) );
AOI21_X1 _17019_ ( .A(fanout_net_38 ), .B1(_03125_ ), .B2(_03128_ ), .ZN(_01089_ ) );
BUF_X8 _17020_ ( .A(_09471_ ), .Z(_03129_ ) );
BUF_X4 _17021_ ( .A(_03129_ ), .Z(_03130_ ) );
NAND4_X1 _17022_ ( .A1(_09994_ ), .A2(_03021_ ), .A3(_03046_ ), .A4(_03130_ ), .ZN(_03131_ ) );
OAI21_X1 _17023_ ( .A(\u_lsu.pmem[5158] ), .B1(_03042_ ), .B2(_03127_ ), .ZN(_03132_ ) );
AOI21_X1 _17024_ ( .A(fanout_net_38 ), .B1(_03131_ ), .B2(_03132_ ), .ZN(_01090_ ) );
BUF_X4 _17025_ ( .A(_03020_ ), .Z(_03133_ ) );
NAND4_X1 _17026_ ( .A1(_09997_ ), .A2(_03133_ ), .A3(_03046_ ), .A4(_03130_ ), .ZN(_03134_ ) );
OAI21_X1 _17027_ ( .A(\u_lsu.pmem[5157] ), .B1(_03042_ ), .B2(_03127_ ), .ZN(_03135_ ) );
AOI21_X1 _17028_ ( .A(fanout_net_39 ), .B1(_03134_ ), .B2(_03135_ ), .ZN(_01091_ ) );
OAI21_X1 _17029_ ( .A(\u_lsu.pmem[5156] ), .B1(_03117_ ), .B2(_03127_ ), .ZN(_03136_ ) );
NAND4_X1 _17030_ ( .A1(_02327_ ), .A2(_03092_ ), .A3(_03112_ ), .A4(_10988_ ), .ZN(_03137_ ) );
AOI21_X1 _17031_ ( .A(fanout_net_39 ), .B1(_03136_ ), .B2(_03137_ ), .ZN(_01092_ ) );
OAI21_X1 _17032_ ( .A(\u_lsu.pmem[5155] ), .B1(_03117_ ), .B2(_03127_ ), .ZN(_03138_ ) );
NAND4_X1 _17033_ ( .A1(_03091_ ), .A2(_03092_ ), .A3(_03112_ ), .A4(_10988_ ), .ZN(_03139_ ) );
AOI21_X1 _17034_ ( .A(fanout_net_39 ), .B1(_03138_ ), .B2(_03139_ ), .ZN(_01093_ ) );
OAI21_X1 _17035_ ( .A(\u_lsu.pmem[5154] ), .B1(_03117_ ), .B2(_03127_ ), .ZN(_03140_ ) );
NAND4_X1 _17036_ ( .A1(_02379_ ), .A2(_03092_ ), .A3(_03112_ ), .A4(_10979_ ), .ZN(_03141_ ) );
AOI21_X1 _17037_ ( .A(fanout_net_39 ), .B1(_03140_ ), .B2(_03141_ ), .ZN(_01094_ ) );
OAI21_X1 _17038_ ( .A(\u_lsu.pmem[5153] ), .B1(_03117_ ), .B2(_03127_ ), .ZN(_03142_ ) );
BUF_X4 _17039_ ( .A(_09616_ ), .Z(_03143_ ) );
NAND4_X1 _17040_ ( .A1(_03143_ ), .A2(_03092_ ), .A3(_03112_ ), .A4(_10979_ ), .ZN(_03144_ ) );
AOI21_X1 _17041_ ( .A(fanout_net_39 ), .B1(_03142_ ), .B2(_03144_ ), .ZN(_01095_ ) );
BUF_X4 _17042_ ( .A(_10015_ ), .Z(_03145_ ) );
NAND2_X1 _17043_ ( .A1(_02996_ ), .A2(_03145_ ), .ZN(_03146_ ) );
OAI21_X1 _17044_ ( .A(\u_lsu.pmem[3650] ), .B1(_02874_ ), .B2(_10501_ ), .ZN(_03147_ ) );
AOI21_X1 _17045_ ( .A(fanout_net_39 ), .B1(_03146_ ), .B2(_03147_ ), .ZN(_01096_ ) );
NAND4_X1 _17046_ ( .A1(_10021_ ), .A2(_03133_ ), .A3(_03046_ ), .A4(_03130_ ), .ZN(_03148_ ) );
OAI21_X1 _17047_ ( .A(\u_lsu.pmem[5152] ), .B1(_03042_ ), .B2(_03127_ ), .ZN(_03149_ ) );
AOI21_X1 _17048_ ( .A(fanout_net_39 ), .B1(_03148_ ), .B2(_03149_ ), .ZN(_01097_ ) );
NAND4_X1 _17049_ ( .A1(_11000_ ), .A2(_10034_ ), .A3(_02500_ ), .A4(_11001_ ), .ZN(_03150_ ) );
AND2_X2 _17050_ ( .A1(_11001_ ), .A2(_09020_ ), .ZN(_03151_ ) );
NAND2_X1 _17051_ ( .A1(_03151_ ), .A2(_10041_ ), .ZN(_03152_ ) );
NAND2_X1 _17052_ ( .A1(_03152_ ), .A2(\u_lsu.pmem[5127] ), .ZN(_03153_ ) );
AOI21_X1 _17053_ ( .A(fanout_net_39 ), .B1(_03150_ ), .B2(_03153_ ), .ZN(_01098_ ) );
INV_X1 _17054_ ( .A(_03151_ ), .ZN(_03154_ ) );
BUF_X2 _17055_ ( .A(_03154_ ), .Z(_03155_ ) );
OR4_X1 _17056_ ( .A1(_09576_ ), .A2(_03155_ ), .A3(_11011_ ), .A4(_10873_ ), .ZN(_03156_ ) );
NAND2_X1 _17057_ ( .A1(_03152_ ), .A2(\u_lsu.pmem[5126] ), .ZN(_03157_ ) );
AOI21_X1 _17058_ ( .A(fanout_net_39 ), .B1(_03156_ ), .B2(_03157_ ), .ZN(_01099_ ) );
OR4_X1 _17059_ ( .A1(_09583_ ), .A2(_03155_ ), .A3(_11011_ ), .A4(_10873_ ), .ZN(_03158_ ) );
NAND2_X1 _17060_ ( .A1(_03152_ ), .A2(\u_lsu.pmem[5125] ), .ZN(_03159_ ) );
AOI21_X1 _17061_ ( .A(fanout_net_39 ), .B1(_03158_ ), .B2(_03159_ ), .ZN(_01100_ ) );
OR4_X1 _17062_ ( .A1(_09146_ ), .A2(_03154_ ), .A3(_02413_ ), .A4(_09498_ ), .ZN(_03160_ ) );
NAND2_X1 _17063_ ( .A1(_03152_ ), .A2(\u_lsu.pmem[5124] ), .ZN(_03161_ ) );
AOI21_X1 _17064_ ( .A(fanout_net_39 ), .B1(_03160_ ), .B2(_03161_ ), .ZN(_01101_ ) );
OR4_X1 _17065_ ( .A1(_09969_ ), .A2(_03154_ ), .A3(_02413_ ), .A4(_09498_ ), .ZN(_03162_ ) );
NAND2_X1 _17066_ ( .A1(_03152_ ), .A2(\u_lsu.pmem[5123] ), .ZN(_03163_ ) );
AOI21_X1 _17067_ ( .A(fanout_net_39 ), .B1(_03162_ ), .B2(_03163_ ), .ZN(_01102_ ) );
NAND4_X1 _17068_ ( .A1(_11021_ ), .A2(_02286_ ), .A3(_03046_ ), .A4(_03130_ ), .ZN(_03164_ ) );
NAND2_X1 _17069_ ( .A1(_03152_ ), .A2(\u_lsu.pmem[5122] ), .ZN(_03165_ ) );
AOI21_X1 _17070_ ( .A(fanout_net_39 ), .B1(_03164_ ), .B2(_03165_ ), .ZN(_01103_ ) );
OR4_X1 _17071_ ( .A1(_09977_ ), .A2(_03154_ ), .A3(_02413_ ), .A4(_09498_ ), .ZN(_03166_ ) );
NAND2_X1 _17072_ ( .A1(_03152_ ), .A2(\u_lsu.pmem[5121] ), .ZN(_03167_ ) );
AOI21_X1 _17073_ ( .A(fanout_net_39 ), .B1(_03166_ ), .B2(_03167_ ), .ZN(_01104_ ) );
OR4_X1 _17074_ ( .A1(_09497_ ), .A2(_03154_ ), .A3(_02413_ ), .A4(_09498_ ), .ZN(_03168_ ) );
NAND2_X1 _17075_ ( .A1(_03152_ ), .A2(\u_lsu.pmem[5120] ), .ZN(_03169_ ) );
AOI21_X1 _17076_ ( .A(fanout_net_39 ), .B1(_03168_ ), .B2(_03169_ ), .ZN(_01105_ ) );
NAND2_X1 _17077_ ( .A1(_02980_ ), .A2(_11030_ ), .ZN(_03170_ ) );
BUF_X4 _17078_ ( .A(_03170_ ), .Z(_03171_ ) );
OAI21_X1 _17079_ ( .A(\u_lsu.pmem[5095] ), .B1(_03117_ ), .B2(_03171_ ), .ZN(_03172_ ) );
NAND4_X1 _17080_ ( .A1(_09742_ ), .A2(_03092_ ), .A3(_03112_ ), .A4(_11030_ ), .ZN(_03173_ ) );
AOI21_X1 _17081_ ( .A(fanout_net_39 ), .B1(_03172_ ), .B2(_03173_ ), .ZN(_01106_ ) );
BUF_X4 _17082_ ( .A(_09616_ ), .Z(_03174_ ) );
NAND2_X1 _17083_ ( .A1(_02996_ ), .A2(_03174_ ), .ZN(_03175_ ) );
OAI21_X1 _17084_ ( .A(\u_lsu.pmem[3649] ), .B1(_02874_ ), .B2(_10501_ ), .ZN(_03176_ ) );
AOI21_X1 _17085_ ( .A(fanout_net_39 ), .B1(_03175_ ), .B2(_03176_ ), .ZN(_01107_ ) );
BUF_X4 _17086_ ( .A(_11453_ ), .Z(_03177_ ) );
NAND4_X1 _17087_ ( .A1(_10062_ ), .A2(_03177_ ), .A3(_03046_ ), .A4(_03130_ ), .ZN(_03178_ ) );
OAI21_X1 _17088_ ( .A(\u_lsu.pmem[5094] ), .B1(_03042_ ), .B2(_03171_ ), .ZN(_03179_ ) );
AOI21_X1 _17089_ ( .A(fanout_net_39 ), .B1(_03178_ ), .B2(_03179_ ), .ZN(_01108_ ) );
NAND4_X1 _17090_ ( .A1(_10075_ ), .A2(_03177_ ), .A3(_03046_ ), .A4(_03130_ ), .ZN(_03180_ ) );
OAI21_X1 _17091_ ( .A(\u_lsu.pmem[5093] ), .B1(_03042_ ), .B2(_03170_ ), .ZN(_03181_ ) );
AOI21_X1 _17092_ ( .A(fanout_net_39 ), .B1(_03180_ ), .B2(_03181_ ), .ZN(_01109_ ) );
NAND4_X1 _17093_ ( .A1(_10079_ ), .A2(_03177_ ), .A3(_03046_ ), .A4(_03130_ ), .ZN(_03182_ ) );
OAI21_X1 _17094_ ( .A(\u_lsu.pmem[5092] ), .B1(_03042_ ), .B2(_03170_ ), .ZN(_03183_ ) );
AOI21_X1 _17095_ ( .A(fanout_net_39 ), .B1(_03182_ ), .B2(_03183_ ), .ZN(_01110_ ) );
NAND4_X1 _17096_ ( .A1(_10084_ ), .A2(_03177_ ), .A3(_03046_ ), .A4(_03130_ ), .ZN(_03184_ ) );
BUF_X4 _17097_ ( .A(_02822_ ), .Z(_03185_ ) );
OAI21_X1 _17098_ ( .A(\u_lsu.pmem[5091] ), .B1(_03185_ ), .B2(_03170_ ), .ZN(_03186_ ) );
AOI21_X1 _17099_ ( .A(fanout_net_39 ), .B1(_03184_ ), .B2(_03186_ ), .ZN(_01111_ ) );
BUF_X4 _17100_ ( .A(_02657_ ), .Z(_03187_ ) );
NAND4_X1 _17101_ ( .A1(_10088_ ), .A2(_03177_ ), .A3(_03187_ ), .A4(_03130_ ), .ZN(_03188_ ) );
OAI21_X1 _17102_ ( .A(\u_lsu.pmem[5090] ), .B1(_03185_ ), .B2(_03170_ ), .ZN(_03189_ ) );
AOI21_X1 _17103_ ( .A(fanout_net_39 ), .B1(_03188_ ), .B2(_03189_ ), .ZN(_01112_ ) );
NAND4_X1 _17104_ ( .A1(_10094_ ), .A2(_03177_ ), .A3(_03187_ ), .A4(_03130_ ), .ZN(_03190_ ) );
OAI21_X1 _17105_ ( .A(\u_lsu.pmem[5089] ), .B1(_03185_ ), .B2(_03170_ ), .ZN(_03191_ ) );
AOI21_X1 _17106_ ( .A(fanout_net_39 ), .B1(_03190_ ), .B2(_03191_ ), .ZN(_01113_ ) );
BUF_X4 _17107_ ( .A(_03129_ ), .Z(_03192_ ) );
NAND4_X1 _17108_ ( .A1(_10098_ ), .A2(_03177_ ), .A3(_03187_ ), .A4(_03192_ ), .ZN(_03193_ ) );
OAI21_X1 _17109_ ( .A(\u_lsu.pmem[5088] ), .B1(_03185_ ), .B2(_03170_ ), .ZN(_03194_ ) );
AOI21_X1 _17110_ ( .A(fanout_net_39 ), .B1(_03193_ ), .B2(_03194_ ), .ZN(_01114_ ) );
NAND2_X1 _17111_ ( .A1(_02980_ ), .A2(_11057_ ), .ZN(_03195_ ) );
BUF_X4 _17112_ ( .A(_03195_ ), .Z(_03196_ ) );
OAI21_X1 _17113_ ( .A(\u_lsu.pmem[5063] ), .B1(_03117_ ), .B2(_03196_ ), .ZN(_03197_ ) );
NAND4_X1 _17114_ ( .A1(_09742_ ), .A2(_03092_ ), .A3(_03112_ ), .A4(_11057_ ), .ZN(_03198_ ) );
AOI21_X1 _17115_ ( .A(fanout_net_39 ), .B1(_03197_ ), .B2(_03198_ ), .ZN(_01115_ ) );
NAND4_X1 _17116_ ( .A1(_10117_ ), .A2(_03177_ ), .A3(_03187_ ), .A4(_03192_ ), .ZN(_03199_ ) );
OAI21_X1 _17117_ ( .A(\u_lsu.pmem[5062] ), .B1(_03185_ ), .B2(_03196_ ), .ZN(_03200_ ) );
AOI21_X1 _17118_ ( .A(fanout_net_39 ), .B1(_03199_ ), .B2(_03200_ ), .ZN(_01116_ ) );
NAND4_X1 _17119_ ( .A1(_10121_ ), .A2(_03177_ ), .A3(_03187_ ), .A4(_03192_ ), .ZN(_03201_ ) );
OAI21_X1 _17120_ ( .A(\u_lsu.pmem[5061] ), .B1(_03185_ ), .B2(_03195_ ), .ZN(_03202_ ) );
AOI21_X1 _17121_ ( .A(fanout_net_39 ), .B1(_03201_ ), .B2(_03202_ ), .ZN(_01117_ ) );
BUF_X4 _17122_ ( .A(_09621_ ), .Z(_03203_ ) );
NAND2_X1 _17123_ ( .A1(_02996_ ), .A2(_03203_ ), .ZN(_03204_ ) );
BUF_X4 _17124_ ( .A(_09562_ ), .Z(_03205_ ) );
OAI21_X1 _17125_ ( .A(\u_lsu.pmem[3648] ), .B1(_03205_ ), .B2(_10501_ ), .ZN(_03206_ ) );
AOI21_X1 _17126_ ( .A(fanout_net_39 ), .B1(_03204_ ), .B2(_03206_ ), .ZN(_01118_ ) );
NAND4_X1 _17127_ ( .A1(_10125_ ), .A2(_03177_ ), .A3(_03187_ ), .A4(_03192_ ), .ZN(_03207_ ) );
OAI21_X1 _17128_ ( .A(\u_lsu.pmem[5060] ), .B1(_03185_ ), .B2(_03195_ ), .ZN(_03208_ ) );
AOI21_X1 _17129_ ( .A(fanout_net_39 ), .B1(_03207_ ), .B2(_03208_ ), .ZN(_01119_ ) );
BUF_X4 _17130_ ( .A(_11453_ ), .Z(_03209_ ) );
NAND4_X1 _17131_ ( .A1(_10131_ ), .A2(_03209_ ), .A3(_03187_ ), .A4(_03192_ ), .ZN(_03210_ ) );
OAI21_X1 _17132_ ( .A(\u_lsu.pmem[5059] ), .B1(_03185_ ), .B2(_03195_ ), .ZN(_03211_ ) );
AOI21_X1 _17133_ ( .A(fanout_net_39 ), .B1(_03210_ ), .B2(_03211_ ), .ZN(_01120_ ) );
NAND4_X1 _17134_ ( .A1(_10135_ ), .A2(_03209_ ), .A3(_03187_ ), .A4(_03192_ ), .ZN(_03212_ ) );
OAI21_X1 _17135_ ( .A(\u_lsu.pmem[5058] ), .B1(_03185_ ), .B2(_03195_ ), .ZN(_03213_ ) );
AOI21_X1 _17136_ ( .A(fanout_net_40 ), .B1(_03212_ ), .B2(_03213_ ), .ZN(_01121_ ) );
NAND4_X1 _17137_ ( .A1(_10138_ ), .A2(_03209_ ), .A3(_03187_ ), .A4(_03192_ ), .ZN(_03214_ ) );
OAI21_X1 _17138_ ( .A(\u_lsu.pmem[5057] ), .B1(_03185_ ), .B2(_03195_ ), .ZN(_03215_ ) );
AOI21_X1 _17139_ ( .A(fanout_net_40 ), .B1(_03214_ ), .B2(_03215_ ), .ZN(_01122_ ) );
NAND4_X1 _17140_ ( .A1(_10144_ ), .A2(_03209_ ), .A3(_03187_ ), .A4(_03192_ ), .ZN(_03216_ ) );
BUF_X4 _17141_ ( .A(_02822_ ), .Z(_03217_ ) );
OAI21_X1 _17142_ ( .A(\u_lsu.pmem[5056] ), .B1(_03217_ ), .B2(_03195_ ), .ZN(_03218_ ) );
AOI21_X1 _17143_ ( .A(fanout_net_40 ), .B1(_03216_ ), .B2(_03218_ ), .ZN(_01123_ ) );
BUF_X4 _17144_ ( .A(_02657_ ), .Z(_03219_ ) );
NAND4_X1 _17145_ ( .A1(_10148_ ), .A2(_03209_ ), .A3(_03219_ ), .A4(_03192_ ), .ZN(_03220_ ) );
NAND2_X1 _17146_ ( .A1(_02980_ ), .A2(_11086_ ), .ZN(_03221_ ) );
BUF_X4 _17147_ ( .A(_03221_ ), .Z(_03222_ ) );
OAI21_X1 _17148_ ( .A(\u_lsu.pmem[5031] ), .B1(_03217_ ), .B2(_03222_ ), .ZN(_03223_ ) );
AOI21_X1 _17149_ ( .A(fanout_net_40 ), .B1(_03220_ ), .B2(_03223_ ), .ZN(_01124_ ) );
NAND4_X1 _17150_ ( .A1(_10156_ ), .A2(_03209_ ), .A3(_03219_ ), .A4(_03192_ ), .ZN(_03224_ ) );
OAI21_X1 _17151_ ( .A(\u_lsu.pmem[5030] ), .B1(_03217_ ), .B2(_03221_ ), .ZN(_03225_ ) );
AOI21_X1 _17152_ ( .A(fanout_net_40 ), .B1(_03224_ ), .B2(_03225_ ), .ZN(_01125_ ) );
BUF_X4 _17153_ ( .A(_03129_ ), .Z(_03226_ ) );
NAND4_X1 _17154_ ( .A1(_10160_ ), .A2(_03209_ ), .A3(_03219_ ), .A4(_03226_ ), .ZN(_03227_ ) );
OAI21_X1 _17155_ ( .A(\u_lsu.pmem[5029] ), .B1(_03217_ ), .B2(_03221_ ), .ZN(_03228_ ) );
AOI21_X1 _17156_ ( .A(fanout_net_40 ), .B1(_03227_ ), .B2(_03228_ ), .ZN(_01126_ ) );
NAND4_X1 _17157_ ( .A1(_10166_ ), .A2(_03209_ ), .A3(_03219_ ), .A4(_03226_ ), .ZN(_03229_ ) );
OAI21_X1 _17158_ ( .A(\u_lsu.pmem[5028] ), .B1(_03217_ ), .B2(_03221_ ), .ZN(_03230_ ) );
AOI21_X1 _17159_ ( .A(fanout_net_40 ), .B1(_03229_ ), .B2(_03230_ ), .ZN(_01127_ ) );
NAND4_X1 _17160_ ( .A1(_10169_ ), .A2(_03209_ ), .A3(_03219_ ), .A4(_03226_ ), .ZN(_03231_ ) );
OAI21_X1 _17161_ ( .A(\u_lsu.pmem[5027] ), .B1(_03217_ ), .B2(_03221_ ), .ZN(_03232_ ) );
AOI21_X1 _17162_ ( .A(fanout_net_40 ), .B1(_03231_ ), .B2(_03232_ ), .ZN(_01128_ ) );
BUF_X4 _17163_ ( .A(_11492_ ), .Z(_03233_ ) );
NAND4_X1 _17164_ ( .A1(_10527_ ), .A2(_03133_ ), .A3(_02429_ ), .A4(_03233_ ), .ZN(_03234_ ) );
OAI21_X1 _17165_ ( .A(\u_lsu.pmem[3623] ), .B1(_03205_ ), .B2(_10533_ ), .ZN(_03235_ ) );
AOI21_X1 _17166_ ( .A(fanout_net_40 ), .B1(_03234_ ), .B2(_03235_ ), .ZN(_01129_ ) );
NAND4_X1 _17167_ ( .A1(_10172_ ), .A2(_03209_ ), .A3(_03219_ ), .A4(_03226_ ), .ZN(_03236_ ) );
OAI21_X1 _17168_ ( .A(\u_lsu.pmem[5026] ), .B1(_03217_ ), .B2(_03221_ ), .ZN(_03237_ ) );
AOI21_X1 _17169_ ( .A(fanout_net_40 ), .B1(_03236_ ), .B2(_03237_ ), .ZN(_01130_ ) );
BUF_X4 _17170_ ( .A(_11453_ ), .Z(_03238_ ) );
NAND4_X1 _17171_ ( .A1(_10176_ ), .A2(_03238_ ), .A3(_03219_ ), .A4(_03226_ ), .ZN(_03239_ ) );
OAI21_X1 _17172_ ( .A(\u_lsu.pmem[5025] ), .B1(_03217_ ), .B2(_03221_ ), .ZN(_03240_ ) );
AOI21_X1 _17173_ ( .A(fanout_net_40 ), .B1(_03239_ ), .B2(_03240_ ), .ZN(_01131_ ) );
OAI21_X1 _17174_ ( .A(\u_lsu.pmem[5024] ), .B1(_03117_ ), .B2(_03222_ ), .ZN(_03241_ ) );
BUF_X4 _17175_ ( .A(_09950_ ), .Z(_03242_ ) );
BUF_X4 _17176_ ( .A(_02881_ ), .Z(_03243_ ) );
NAND4_X1 _17177_ ( .A1(_02720_ ), .A2(_03242_ ), .A3(_03243_ ), .A4(_11086_ ), .ZN(_03244_ ) );
AOI21_X1 _17178_ ( .A(fanout_net_40 ), .B1(_03241_ ), .B2(_03244_ ), .ZN(_01132_ ) );
NAND2_X1 _17179_ ( .A1(_11108_ ), .A2(_09475_ ), .ZN(_03245_ ) );
BUF_X4 _17180_ ( .A(_03245_ ), .Z(_03246_ ) );
OAI21_X1 _17181_ ( .A(\u_lsu.pmem[4999] ), .B1(_03246_ ), .B2(_03070_ ), .ZN(_03247_ ) );
NAND4_X1 _17182_ ( .A1(_11113_ ), .A2(_10752_ ), .A3(_03243_ ), .A4(_03119_ ), .ZN(_03248_ ) );
AOI21_X1 _17183_ ( .A(fanout_net_40 ), .B1(_03247_ ), .B2(_03248_ ), .ZN(_01133_ ) );
OAI21_X1 _17184_ ( .A(\u_lsu.pmem[4998] ), .B1(_03246_ ), .B2(_03070_ ), .ZN(_03249_ ) );
NAND4_X1 _17185_ ( .A1(_11113_ ), .A2(_03056_ ), .A3(_03243_ ), .A4(_03119_ ), .ZN(_03250_ ) );
AOI21_X1 _17186_ ( .A(fanout_net_40 ), .B1(_03249_ ), .B2(_03250_ ), .ZN(_01134_ ) );
OAI21_X1 _17187_ ( .A(\u_lsu.pmem[4997] ), .B1(_03246_ ), .B2(_03070_ ), .ZN(_03251_ ) );
NAND4_X1 _17188_ ( .A1(_11113_ ), .A2(_03059_ ), .A3(_03243_ ), .A4(_03119_ ), .ZN(_03252_ ) );
AOI21_X1 _17189_ ( .A(fanout_net_40 ), .B1(_03251_ ), .B2(_03252_ ), .ZN(_01135_ ) );
OAI21_X1 _17190_ ( .A(\u_lsu.pmem[4996] ), .B1(_03246_ ), .B2(_03070_ ), .ZN(_03253_ ) );
BUF_X4 _17191_ ( .A(_11112_ ), .Z(_03254_ ) );
NAND4_X1 _17192_ ( .A1(_03254_ ), .A2(_03064_ ), .A3(_03243_ ), .A4(_03119_ ), .ZN(_03255_ ) );
AOI21_X1 _17193_ ( .A(fanout_net_40 ), .B1(_03253_ ), .B2(_03255_ ), .ZN(_01136_ ) );
OAI21_X1 _17194_ ( .A(\u_lsu.pmem[4995] ), .B1(_03246_ ), .B2(_03070_ ), .ZN(_03256_ ) );
NAND4_X1 _17195_ ( .A1(_03254_ ), .A2(_10915_ ), .A3(_03243_ ), .A4(_03119_ ), .ZN(_03257_ ) );
AOI21_X1 _17196_ ( .A(fanout_net_40 ), .B1(_03256_ ), .B2(_03257_ ), .ZN(_01137_ ) );
OAI21_X1 _17197_ ( .A(\u_lsu.pmem[4994] ), .B1(_03246_ ), .B2(_03070_ ), .ZN(_03258_ ) );
NAND4_X1 _17198_ ( .A1(_09874_ ), .A2(_11536_ ), .A3(_03243_ ), .A4(_03119_ ), .ZN(_03259_ ) );
AOI21_X1 _17199_ ( .A(fanout_net_40 ), .B1(_03258_ ), .B2(_03259_ ), .ZN(_01138_ ) );
OAI21_X1 _17200_ ( .A(\u_lsu.pmem[4993] ), .B1(_03246_ ), .B2(_03070_ ), .ZN(_03260_ ) );
NAND4_X1 _17201_ ( .A1(_03254_ ), .A2(_02308_ ), .A3(_03243_ ), .A4(_03119_ ), .ZN(_03261_ ) );
AOI21_X1 _17202_ ( .A(fanout_net_40 ), .B1(_03260_ ), .B2(_03261_ ), .ZN(_01139_ ) );
NAND4_X1 _17203_ ( .A1(_09787_ ), .A2(_03238_ ), .A3(_03219_ ), .A4(_03226_ ), .ZN(_03262_ ) );
OAI21_X1 _17204_ ( .A(\u_lsu.pmem[4321] ), .B1(_03217_ ), .B2(_09751_ ), .ZN(_03263_ ) );
AOI21_X1 _17205_ ( .A(fanout_net_40 ), .B1(_03262_ ), .B2(_03263_ ), .ZN(_01140_ ) );
NAND4_X1 _17206_ ( .A1(_10535_ ), .A2(_03133_ ), .A3(_02429_ ), .A4(_03233_ ), .ZN(_03264_ ) );
OAI21_X1 _17207_ ( .A(\u_lsu.pmem[3622] ), .B1(_03205_ ), .B2(_10533_ ), .ZN(_03265_ ) );
AOI21_X1 _17208_ ( .A(fanout_net_40 ), .B1(_03264_ ), .B2(_03265_ ), .ZN(_01141_ ) );
OAI21_X1 _17209_ ( .A(\u_lsu.pmem[4992] ), .B1(_03246_ ), .B2(_03070_ ), .ZN(_03266_ ) );
BUF_X4 _17210_ ( .A(_10904_ ), .Z(_03267_ ) );
NAND4_X1 _17211_ ( .A1(_03254_ ), .A2(_11131_ ), .A3(_03243_ ), .A4(_03267_ ), .ZN(_03268_ ) );
AOI21_X1 _17212_ ( .A(fanout_net_40 ), .B1(_03266_ ), .B2(_03268_ ), .ZN(_01142_ ) );
BUF_X4 _17213_ ( .A(_09459_ ), .Z(_03269_ ) );
INV_X1 _17214_ ( .A(_11133_ ), .ZN(_03270_ ) );
NOR2_X1 _17215_ ( .A1(_09134_ ), .A2(_03270_ ), .ZN(_03271_ ) );
INV_X1 _17216_ ( .A(_03271_ ), .ZN(_03272_ ) );
BUF_X4 _17217_ ( .A(_03272_ ), .Z(_03273_ ) );
OAI21_X1 _17218_ ( .A(\u_lsu.pmem[4967] ), .B1(_03269_ ), .B2(_03273_ ), .ZN(_03274_ ) );
BUF_X4 _17219_ ( .A(_09635_ ), .Z(_03275_ ) );
BUF_X4 _17220_ ( .A(_03271_ ), .Z(_03276_ ) );
NAND3_X1 _17221_ ( .A1(_11000_ ), .A2(_03275_ ), .A3(_03276_ ), .ZN(_03277_ ) );
AOI21_X1 _17222_ ( .A(fanout_net_40 ), .B1(_03274_ ), .B2(_03277_ ), .ZN(_01143_ ) );
OAI21_X1 _17223_ ( .A(\u_lsu.pmem[4966] ), .B1(_03269_ ), .B2(_03273_ ), .ZN(_03278_ ) );
NAND3_X1 _17224_ ( .A1(_10719_ ), .A2(_03275_ ), .A3(_03276_ ), .ZN(_03279_ ) );
AOI21_X1 _17225_ ( .A(fanout_net_40 ), .B1(_03278_ ), .B2(_03279_ ), .ZN(_01144_ ) );
OAI21_X1 _17226_ ( .A(\u_lsu.pmem[4965] ), .B1(_03269_ ), .B2(_03272_ ), .ZN(_03280_ ) );
NAND3_X1 _17227_ ( .A1(_10728_ ), .A2(_03275_ ), .A3(_03271_ ), .ZN(_03281_ ) );
AOI21_X1 _17228_ ( .A(fanout_net_40 ), .B1(_03280_ ), .B2(_03281_ ), .ZN(_01145_ ) );
OAI21_X1 _17229_ ( .A(\u_lsu.pmem[4964] ), .B1(_03269_ ), .B2(_03272_ ), .ZN(_03282_ ) );
NAND3_X1 _17230_ ( .A1(_11152_ ), .A2(_03275_ ), .A3(_03271_ ), .ZN(_03283_ ) );
AOI21_X1 _17231_ ( .A(fanout_net_40 ), .B1(_03282_ ), .B2(_03283_ ), .ZN(_01146_ ) );
OAI21_X1 _17232_ ( .A(\u_lsu.pmem[4963] ), .B1(_03269_ ), .B2(_03272_ ), .ZN(_03284_ ) );
NAND3_X1 _17233_ ( .A1(_10733_ ), .A2(_03275_ ), .A3(_03271_ ), .ZN(_03285_ ) );
AOI21_X1 _17234_ ( .A(fanout_net_40 ), .B1(_03284_ ), .B2(_03285_ ), .ZN(_01147_ ) );
OAI21_X1 _17235_ ( .A(\u_lsu.pmem[4962] ), .B1(_03269_ ), .B2(_03272_ ), .ZN(_03286_ ) );
NAND3_X1 _17236_ ( .A1(_11158_ ), .A2(_03275_ ), .A3(_03271_ ), .ZN(_03287_ ) );
AOI21_X1 _17237_ ( .A(fanout_net_40 ), .B1(_03286_ ), .B2(_03287_ ), .ZN(_01148_ ) );
OAI21_X1 _17238_ ( .A(\u_lsu.pmem[4961] ), .B1(_03269_ ), .B2(_03272_ ), .ZN(_03288_ ) );
NAND3_X1 _17239_ ( .A1(_10738_ ), .A2(_03275_ ), .A3(_03271_ ), .ZN(_03289_ ) );
AOI21_X1 _17240_ ( .A(fanout_net_40 ), .B1(_03288_ ), .B2(_03289_ ), .ZN(_01149_ ) );
OAI21_X1 _17241_ ( .A(\u_lsu.pmem[4960] ), .B1(_03269_ ), .B2(_03272_ ), .ZN(_03290_ ) );
NAND3_X1 _17242_ ( .A1(_10741_ ), .A2(_03275_ ), .A3(_03271_ ), .ZN(_03291_ ) );
AOI21_X1 _17243_ ( .A(fanout_net_40 ), .B1(_03290_ ), .B2(_03291_ ), .ZN(_01150_ ) );
INV_X1 _17244_ ( .A(_11168_ ), .ZN(_03292_ ) );
NOR2_X1 _17245_ ( .A1(_09134_ ), .A2(_03292_ ), .ZN(_03293_ ) );
INV_X1 _17246_ ( .A(_03293_ ), .ZN(_03294_ ) );
BUF_X4 _17247_ ( .A(_03294_ ), .Z(_03295_ ) );
OAI21_X1 _17248_ ( .A(\u_lsu.pmem[4935] ), .B1(_03269_ ), .B2(_03295_ ), .ZN(_03296_ ) );
BUF_X4 _17249_ ( .A(_03293_ ), .Z(_03297_ ) );
NAND3_X1 _17250_ ( .A1(_11000_ ), .A2(_03275_ ), .A3(_03297_ ), .ZN(_03298_ ) );
AOI21_X1 _17251_ ( .A(fanout_net_41 ), .B1(_03296_ ), .B2(_03298_ ), .ZN(_01151_ ) );
BUF_X4 _17252_ ( .A(_02196_ ), .Z(_03299_ ) );
NAND4_X1 _17253_ ( .A1(_10538_ ), .A2(_03133_ ), .A3(_03299_ ), .A4(_03233_ ), .ZN(_03300_ ) );
OAI21_X1 _17254_ ( .A(\u_lsu.pmem[3621] ), .B1(_03205_ ), .B2(_10532_ ), .ZN(_03301_ ) );
AOI21_X1 _17255_ ( .A(fanout_net_41 ), .B1(_03300_ ), .B2(_03301_ ), .ZN(_01152_ ) );
OAI21_X1 _17256_ ( .A(\u_lsu.pmem[4934] ), .B1(_03269_ ), .B2(_03295_ ), .ZN(_03302_ ) );
NAND3_X1 _17257_ ( .A1(_10719_ ), .A2(_03275_ ), .A3(_03297_ ), .ZN(_03303_ ) );
AOI21_X1 _17258_ ( .A(fanout_net_41 ), .B1(_03302_ ), .B2(_03303_ ), .ZN(_01153_ ) );
BUF_X4 _17259_ ( .A(_09459_ ), .Z(_03304_ ) );
OAI21_X1 _17260_ ( .A(\u_lsu.pmem[4933] ), .B1(_03304_ ), .B2(_03294_ ), .ZN(_03305_ ) );
BUF_X4 _17261_ ( .A(_09635_ ), .Z(_03306_ ) );
NAND3_X1 _17262_ ( .A1(_10728_ ), .A2(_03306_ ), .A3(_03293_ ), .ZN(_03307_ ) );
AOI21_X1 _17263_ ( .A(fanout_net_41 ), .B1(_03305_ ), .B2(_03307_ ), .ZN(_01154_ ) );
OAI21_X1 _17264_ ( .A(\u_lsu.pmem[4932] ), .B1(_03304_ ), .B2(_03294_ ), .ZN(_03308_ ) );
NAND3_X1 _17265_ ( .A1(_11152_ ), .A2(_03306_ ), .A3(_03293_ ), .ZN(_03309_ ) );
AOI21_X1 _17266_ ( .A(fanout_net_41 ), .B1(_03308_ ), .B2(_03309_ ), .ZN(_01155_ ) );
OAI21_X1 _17267_ ( .A(\u_lsu.pmem[4931] ), .B1(_03304_ ), .B2(_03294_ ), .ZN(_03310_ ) );
NAND3_X1 _17268_ ( .A1(_10733_ ), .A2(_03306_ ), .A3(_03293_ ), .ZN(_03311_ ) );
AOI21_X1 _17269_ ( .A(fanout_net_41 ), .B1(_03310_ ), .B2(_03311_ ), .ZN(_01156_ ) );
OAI21_X1 _17270_ ( .A(\u_lsu.pmem[4930] ), .B1(_03304_ ), .B2(_03294_ ), .ZN(_03312_ ) );
NAND3_X1 _17271_ ( .A1(_09612_ ), .A2(_03306_ ), .A3(_03293_ ), .ZN(_03313_ ) );
AOI21_X1 _17272_ ( .A(fanout_net_41 ), .B1(_03312_ ), .B2(_03313_ ), .ZN(_01157_ ) );
OAI21_X1 _17273_ ( .A(\u_lsu.pmem[4929] ), .B1(_03304_ ), .B2(_03294_ ), .ZN(_03314_ ) );
NAND3_X1 _17274_ ( .A1(_10738_ ), .A2(_03306_ ), .A3(_03293_ ), .ZN(_03315_ ) );
AOI21_X1 _17275_ ( .A(fanout_net_41 ), .B1(_03314_ ), .B2(_03315_ ), .ZN(_01158_ ) );
OAI21_X1 _17276_ ( .A(\u_lsu.pmem[4928] ), .B1(_03304_ ), .B2(_03294_ ), .ZN(_03316_ ) );
NAND3_X1 _17277_ ( .A1(_10741_ ), .A2(_03306_ ), .A3(_03293_ ), .ZN(_03317_ ) );
AOI21_X1 _17278_ ( .A(fanout_net_41 ), .B1(_03316_ ), .B2(_03317_ ), .ZN(_01159_ ) );
NAND4_X1 _17279_ ( .A1(_10250_ ), .A2(_03238_ ), .A3(_03219_ ), .A4(_03226_ ), .ZN(_03318_ ) );
INV_X1 _17280_ ( .A(_11197_ ), .ZN(_03319_ ) );
NOR2_X4 _17281_ ( .A1(_10325_ ), .A2(_03319_ ), .ZN(_03320_ ) );
INV_X1 _17282_ ( .A(_03320_ ), .ZN(_03321_ ) );
OAI21_X1 _17283_ ( .A(\u_lsu.pmem[4903] ), .B1(_03217_ ), .B2(_03321_ ), .ZN(_03322_ ) );
AOI21_X1 _17284_ ( .A(fanout_net_41 ), .B1(_03318_ ), .B2(_03322_ ), .ZN(_01160_ ) );
NAND4_X1 _17285_ ( .A1(_10263_ ), .A2(_03238_ ), .A3(_03219_ ), .A4(_03226_ ), .ZN(_03323_ ) );
BUF_X4 _17286_ ( .A(_02822_ ), .Z(_03324_ ) );
OAI21_X1 _17287_ ( .A(\u_lsu.pmem[4902] ), .B1(_03324_ ), .B2(_03321_ ), .ZN(_03325_ ) );
AOI21_X1 _17288_ ( .A(fanout_net_41 ), .B1(_03323_ ), .B2(_03325_ ), .ZN(_01161_ ) );
BUF_X8 _17289_ ( .A(_09455_ ), .Z(_03326_ ) );
BUF_X4 _17290_ ( .A(_03326_ ), .Z(_03327_ ) );
NAND4_X1 _17291_ ( .A1(_10267_ ), .A2(_03238_ ), .A3(_03327_ ), .A4(_03226_ ), .ZN(_03328_ ) );
OAI21_X1 _17292_ ( .A(\u_lsu.pmem[4901] ), .B1(_03324_ ), .B2(_03321_ ), .ZN(_03329_ ) );
AOI21_X1 _17293_ ( .A(fanout_net_41 ), .B1(_03328_ ), .B2(_03329_ ), .ZN(_01162_ ) );
NOR2_X1 _17294_ ( .A1(_11159_ ), .A2(_10532_ ), .ZN(_03330_ ) );
NAND2_X1 _17295_ ( .A1(_03330_ ), .A2(_03084_ ), .ZN(_03331_ ) );
OAI21_X1 _17296_ ( .A(\u_lsu.pmem[3620] ), .B1(_03205_ ), .B2(_10532_ ), .ZN(_03332_ ) );
AOI21_X1 _17297_ ( .A(fanout_net_41 ), .B1(_03331_ ), .B2(_03332_ ), .ZN(_01163_ ) );
AND2_X1 _17298_ ( .A1(_09141_ ), .A2(_03320_ ), .ZN(_03333_ ) );
OAI21_X1 _17299_ ( .A(_10715_ ), .B1(_03333_ ), .B2(\u_lsu.pmem[4900] ), .ZN(_03334_ ) );
AOI21_X1 _17300_ ( .A(_03334_ ), .B1(_09691_ ), .B2(_03333_ ), .ZN(_01164_ ) );
BUF_X4 _17301_ ( .A(_03321_ ), .Z(_03335_ ) );
OAI21_X1 _17302_ ( .A(\u_lsu.pmem[4899] ), .B1(_03304_ ), .B2(_03335_ ), .ZN(_03336_ ) );
NAND3_X1 _17303_ ( .A1(_10733_ ), .A2(_03306_ ), .A3(_03320_ ), .ZN(_03337_ ) );
AOI21_X1 _17304_ ( .A(fanout_net_41 ), .B1(_03336_ ), .B2(_03337_ ), .ZN(_01165_ ) );
OAI21_X1 _17305_ ( .A(\u_lsu.pmem[4898] ), .B1(_03304_ ), .B2(_03335_ ), .ZN(_03338_ ) );
NAND3_X1 _17306_ ( .A1(_09612_ ), .A2(_03306_ ), .A3(_03320_ ), .ZN(_03339_ ) );
AOI21_X1 _17307_ ( .A(fanout_net_41 ), .B1(_03338_ ), .B2(_03339_ ), .ZN(_01166_ ) );
OAI21_X1 _17308_ ( .A(\u_lsu.pmem[4897] ), .B1(_03304_ ), .B2(_03335_ ), .ZN(_03340_ ) );
NAND3_X1 _17309_ ( .A1(_10738_ ), .A2(_03306_ ), .A3(_03320_ ), .ZN(_03341_ ) );
AOI21_X1 _17310_ ( .A(fanout_net_41 ), .B1(_03340_ ), .B2(_03341_ ), .ZN(_01167_ ) );
NAND4_X1 _17311_ ( .A1(_10279_ ), .A2(_03238_ ), .A3(_03327_ ), .A4(_03226_ ), .ZN(_03342_ ) );
OAI21_X1 _17312_ ( .A(\u_lsu.pmem[4896] ), .B1(_03324_ ), .B2(_03321_ ), .ZN(_03343_ ) );
AOI21_X1 _17313_ ( .A(fanout_net_41 ), .B1(_03342_ ), .B2(_03343_ ), .ZN(_01168_ ) );
BUF_X4 _17314_ ( .A(_03129_ ), .Z(_03344_ ) );
NAND4_X1 _17315_ ( .A1(_10285_ ), .A2(_03238_ ), .A3(_03327_ ), .A4(_03344_ ), .ZN(_03345_ ) );
NAND3_X1 _17316_ ( .A1(_09454_ ), .A2(_09842_ ), .A3(_10289_ ), .ZN(_03346_ ) );
BUF_X4 _17317_ ( .A(_03346_ ), .Z(_03347_ ) );
OAI21_X1 _17318_ ( .A(\u_lsu.pmem[4871] ), .B1(_03324_ ), .B2(_03347_ ), .ZN(_03348_ ) );
AOI21_X1 _17319_ ( .A(fanout_net_41 ), .B1(_03345_ ), .B2(_03348_ ), .ZN(_01169_ ) );
NAND4_X1 _17320_ ( .A1(_10295_ ), .A2(_03238_ ), .A3(_03327_ ), .A4(_03344_ ), .ZN(_03349_ ) );
OAI21_X1 _17321_ ( .A(\u_lsu.pmem[4870] ), .B1(_03324_ ), .B2(_03346_ ), .ZN(_03350_ ) );
AOI21_X1 _17322_ ( .A(fanout_net_41 ), .B1(_03349_ ), .B2(_03350_ ), .ZN(_01170_ ) );
NAND4_X1 _17323_ ( .A1(_10299_ ), .A2(_03238_ ), .A3(_03327_ ), .A4(_03344_ ), .ZN(_03351_ ) );
OAI21_X1 _17324_ ( .A(\u_lsu.pmem[4869] ), .B1(_03324_ ), .B2(_03346_ ), .ZN(_03352_ ) );
AOI21_X1 _17325_ ( .A(fanout_net_41 ), .B1(_03351_ ), .B2(_03352_ ), .ZN(_01171_ ) );
NAND4_X1 _17326_ ( .A1(_10306_ ), .A2(_03238_ ), .A3(_03327_ ), .A4(_03344_ ), .ZN(_03353_ ) );
OAI21_X1 _17327_ ( .A(\u_lsu.pmem[4868] ), .B1(_03324_ ), .B2(_03346_ ), .ZN(_03354_ ) );
AOI21_X1 _17328_ ( .A(fanout_net_41 ), .B1(_03353_ ), .B2(_03354_ ), .ZN(_01172_ ) );
BUF_X4 _17329_ ( .A(_11453_ ), .Z(_03355_ ) );
NAND4_X1 _17330_ ( .A1(_10309_ ), .A2(_03355_ ), .A3(_03327_ ), .A4(_03344_ ), .ZN(_03356_ ) );
OAI21_X1 _17331_ ( .A(\u_lsu.pmem[4867] ), .B1(_03324_ ), .B2(_03346_ ), .ZN(_03357_ ) );
AOI21_X1 _17332_ ( .A(fanout_net_41 ), .B1(_03356_ ), .B2(_03357_ ), .ZN(_01173_ ) );
NAND2_X1 _17333_ ( .A1(_03330_ ), .A2(_03114_ ), .ZN(_03358_ ) );
OAI21_X1 _17334_ ( .A(\u_lsu.pmem[3619] ), .B1(_03205_ ), .B2(_10532_ ), .ZN(_03359_ ) );
AOI21_X1 _17335_ ( .A(fanout_net_41 ), .B1(_03358_ ), .B2(_03359_ ), .ZN(_01174_ ) );
OAI21_X1 _17336_ ( .A(\u_lsu.pmem[4866] ), .B1(_03304_ ), .B2(_03347_ ), .ZN(_03360_ ) );
BUF_X4 _17337_ ( .A(_09883_ ), .Z(_03361_ ) );
NAND4_X1 _17338_ ( .A1(_09510_ ), .A2(_03361_ ), .A3(_03243_ ), .A4(_10313_ ), .ZN(_03362_ ) );
AOI21_X1 _17339_ ( .A(fanout_net_41 ), .B1(_03360_ ), .B2(_03362_ ), .ZN(_01175_ ) );
NAND4_X1 _17340_ ( .A1(_10316_ ), .A2(_03355_ ), .A3(_03327_ ), .A4(_03344_ ), .ZN(_03363_ ) );
OAI21_X1 _17341_ ( .A(\u_lsu.pmem[4865] ), .B1(_03324_ ), .B2(_03346_ ), .ZN(_03364_ ) );
AOI21_X1 _17342_ ( .A(fanout_net_41 ), .B1(_03363_ ), .B2(_03364_ ), .ZN(_01176_ ) );
NAND4_X1 _17343_ ( .A1(_10320_ ), .A2(_03355_ ), .A3(_03327_ ), .A4(_03344_ ), .ZN(_03365_ ) );
OAI21_X1 _17344_ ( .A(\u_lsu.pmem[4864] ), .B1(_03324_ ), .B2(_03346_ ), .ZN(_03366_ ) );
AOI21_X1 _17345_ ( .A(fanout_net_41 ), .B1(_03365_ ), .B2(_03366_ ), .ZN(_01177_ ) );
BUF_X4 _17346_ ( .A(_09459_ ), .Z(_03367_ ) );
NAND2_X1 _17347_ ( .A1(_02980_ ), .A2(_11245_ ), .ZN(_03368_ ) );
BUF_X4 _17348_ ( .A(_03368_ ), .Z(_03369_ ) );
OAI21_X1 _17349_ ( .A(\u_lsu.pmem[4839] ), .B1(_03367_ ), .B2(_03369_ ), .ZN(_03370_ ) );
BUF_X4 _17350_ ( .A(_02881_ ), .Z(_03371_ ) );
NAND4_X1 _17351_ ( .A1(_09742_ ), .A2(_03242_ ), .A3(_03371_ ), .A4(_11245_ ), .ZN(_03372_ ) );
AOI21_X1 _17352_ ( .A(fanout_net_41 ), .B1(_03370_ ), .B2(_03372_ ), .ZN(_01178_ ) );
NAND4_X1 _17353_ ( .A1(_10332_ ), .A2(_03355_ ), .A3(_03327_ ), .A4(_03344_ ), .ZN(_03373_ ) );
BUF_X4 _17354_ ( .A(_02822_ ), .Z(_03374_ ) );
OAI21_X1 _17355_ ( .A(\u_lsu.pmem[4838] ), .B1(_03374_ ), .B2(_03369_ ), .ZN(_03375_ ) );
AOI21_X1 _17356_ ( .A(fanout_net_41 ), .B1(_03373_ ), .B2(_03375_ ), .ZN(_01179_ ) );
BUF_X4 _17357_ ( .A(_03326_ ), .Z(_03376_ ) );
NAND4_X1 _17358_ ( .A1(_10336_ ), .A2(_03355_ ), .A3(_03376_ ), .A4(_03344_ ), .ZN(_03377_ ) );
OAI21_X1 _17359_ ( .A(\u_lsu.pmem[4837] ), .B1(_03374_ ), .B2(_03368_ ), .ZN(_03378_ ) );
AOI21_X1 _17360_ ( .A(fanout_net_41 ), .B1(_03377_ ), .B2(_03378_ ), .ZN(_01180_ ) );
NAND4_X1 _17361_ ( .A1(_10339_ ), .A2(_03355_ ), .A3(_03376_ ), .A4(_03344_ ), .ZN(_03379_ ) );
OAI21_X1 _17362_ ( .A(\u_lsu.pmem[4836] ), .B1(_03374_ ), .B2(_03368_ ), .ZN(_03380_ ) );
AOI21_X1 _17363_ ( .A(fanout_net_41 ), .B1(_03379_ ), .B2(_03380_ ), .ZN(_01181_ ) );
BUF_X4 _17364_ ( .A(_03129_ ), .Z(_03381_ ) );
NAND4_X1 _17365_ ( .A1(_10345_ ), .A2(_03355_ ), .A3(_03376_ ), .A4(_03381_ ), .ZN(_03382_ ) );
OAI21_X1 _17366_ ( .A(\u_lsu.pmem[4835] ), .B1(_03374_ ), .B2(_03368_ ), .ZN(_03383_ ) );
AOI21_X1 _17367_ ( .A(fanout_net_42 ), .B1(_03382_ ), .B2(_03383_ ), .ZN(_01182_ ) );
NAND4_X1 _17368_ ( .A1(_10350_ ), .A2(_03355_ ), .A3(_03376_ ), .A4(_03381_ ), .ZN(_03384_ ) );
OAI21_X1 _17369_ ( .A(\u_lsu.pmem[4834] ), .B1(_03374_ ), .B2(_03368_ ), .ZN(_03385_ ) );
AOI21_X1 _17370_ ( .A(fanout_net_42 ), .B1(_03384_ ), .B2(_03385_ ), .ZN(_01183_ ) );
NAND4_X1 _17371_ ( .A1(_10354_ ), .A2(_03355_ ), .A3(_03376_ ), .A4(_03381_ ), .ZN(_03386_ ) );
OAI21_X1 _17372_ ( .A(\u_lsu.pmem[4833] ), .B1(_03374_ ), .B2(_03368_ ), .ZN(_03387_ ) );
AOI21_X1 _17373_ ( .A(fanout_net_42 ), .B1(_03386_ ), .B2(_03387_ ), .ZN(_01184_ ) );
NAND2_X1 _17374_ ( .A1(_03330_ ), .A2(_03145_ ), .ZN(_03388_ ) );
OAI21_X1 _17375_ ( .A(\u_lsu.pmem[3618] ), .B1(_03205_ ), .B2(_10532_ ), .ZN(_03389_ ) );
AOI21_X1 _17376_ ( .A(fanout_net_42 ), .B1(_03388_ ), .B2(_03389_ ), .ZN(_01185_ ) );
NAND4_X1 _17377_ ( .A1(_10357_ ), .A2(_03355_ ), .A3(_03376_ ), .A4(_03381_ ), .ZN(_03390_ ) );
OAI21_X1 _17378_ ( .A(\u_lsu.pmem[4832] ), .B1(_03374_ ), .B2(_03368_ ), .ZN(_03391_ ) );
AOI21_X1 _17379_ ( .A(fanout_net_42 ), .B1(_03390_ ), .B2(_03391_ ), .ZN(_01186_ ) );
NAND2_X1 _17380_ ( .A1(_02980_ ), .A2(_11267_ ), .ZN(_03392_ ) );
BUF_X4 _17381_ ( .A(_03392_ ), .Z(_03393_ ) );
OAI21_X1 _17382_ ( .A(\u_lsu.pmem[4807] ), .B1(_03367_ ), .B2(_03393_ ), .ZN(_03394_ ) );
NAND4_X1 _17383_ ( .A1(_09742_ ), .A2(_03242_ ), .A3(_03371_ ), .A4(_11267_ ), .ZN(_03395_ ) );
AOI21_X1 _17384_ ( .A(fanout_net_42 ), .B1(_03394_ ), .B2(_03395_ ), .ZN(_01187_ ) );
BUF_X8 _17385_ ( .A(_09539_ ), .Z(_03396_ ) );
BUF_X4 _17386_ ( .A(_03396_ ), .Z(_03397_ ) );
NAND4_X1 _17387_ ( .A1(_10368_ ), .A2(_03397_ ), .A3(_03376_ ), .A4(_03381_ ), .ZN(_03398_ ) );
OAI21_X1 _17388_ ( .A(\u_lsu.pmem[4806] ), .B1(_03374_ ), .B2(_03393_ ), .ZN(_03399_ ) );
AOI21_X1 _17389_ ( .A(fanout_net_42 ), .B1(_03398_ ), .B2(_03399_ ), .ZN(_01188_ ) );
NAND4_X1 _17390_ ( .A1(_10371_ ), .A2(_03397_ ), .A3(_03376_ ), .A4(_03381_ ), .ZN(_03400_ ) );
OAI21_X1 _17391_ ( .A(\u_lsu.pmem[4805] ), .B1(_03374_ ), .B2(_03392_ ), .ZN(_03401_ ) );
AOI21_X1 _17392_ ( .A(fanout_net_42 ), .B1(_03400_ ), .B2(_03401_ ), .ZN(_01189_ ) );
NAND4_X1 _17393_ ( .A1(_10374_ ), .A2(_03397_ ), .A3(_03376_ ), .A4(_03381_ ), .ZN(_03402_ ) );
OAI21_X1 _17394_ ( .A(\u_lsu.pmem[4804] ), .B1(_03374_ ), .B2(_03392_ ), .ZN(_03403_ ) );
AOI21_X1 _17395_ ( .A(fanout_net_42 ), .B1(_03402_ ), .B2(_03403_ ), .ZN(_01190_ ) );
NAND4_X1 _17396_ ( .A1(_10377_ ), .A2(_03397_ ), .A3(_03376_ ), .A4(_03381_ ), .ZN(_03404_ ) );
BUF_X4 _17397_ ( .A(_02822_ ), .Z(_03405_ ) );
OAI21_X1 _17398_ ( .A(\u_lsu.pmem[4803] ), .B1(_03405_ ), .B2(_03392_ ), .ZN(_03406_ ) );
AOI21_X1 _17399_ ( .A(fanout_net_42 ), .B1(_03404_ ), .B2(_03406_ ), .ZN(_01191_ ) );
BUF_X4 _17400_ ( .A(_03326_ ), .Z(_03407_ ) );
NAND4_X1 _17401_ ( .A1(_10381_ ), .A2(_03397_ ), .A3(_03407_ ), .A4(_03381_ ), .ZN(_03408_ ) );
OAI21_X1 _17402_ ( .A(\u_lsu.pmem[4802] ), .B1(_03405_ ), .B2(_03392_ ), .ZN(_03409_ ) );
AOI21_X1 _17403_ ( .A(fanout_net_42 ), .B1(_03408_ ), .B2(_03409_ ), .ZN(_01192_ ) );
NAND4_X1 _17404_ ( .A1(_10384_ ), .A2(_03397_ ), .A3(_03407_ ), .A4(_03381_ ), .ZN(_03410_ ) );
OAI21_X1 _17405_ ( .A(\u_lsu.pmem[4801] ), .B1(_03405_ ), .B2(_03392_ ), .ZN(_03411_ ) );
AOI21_X1 _17406_ ( .A(fanout_net_42 ), .B1(_03410_ ), .B2(_03411_ ), .ZN(_01193_ ) );
BUF_X4 _17407_ ( .A(_03129_ ), .Z(_03412_ ) );
NAND4_X1 _17408_ ( .A1(_10391_ ), .A2(_03397_ ), .A3(_03407_ ), .A4(_03412_ ), .ZN(_03413_ ) );
OAI21_X1 _17409_ ( .A(\u_lsu.pmem[4800] ), .B1(_03405_ ), .B2(_03392_ ), .ZN(_03414_ ) );
AOI21_X1 _17410_ ( .A(fanout_net_42 ), .B1(_03413_ ), .B2(_03414_ ), .ZN(_01194_ ) );
NAND4_X1 _17411_ ( .A1(_10394_ ), .A2(_03397_ ), .A3(_03407_ ), .A4(_03412_ ), .ZN(_03415_ ) );
NAND2_X1 _17412_ ( .A1(_11292_ ), .A2(_02484_ ), .ZN(_03416_ ) );
BUF_X4 _17413_ ( .A(_03416_ ), .Z(_03417_ ) );
OAI21_X1 _17414_ ( .A(\u_lsu.pmem[4775] ), .B1(_03405_ ), .B2(_03417_ ), .ZN(_03418_ ) );
AOI21_X1 _17415_ ( .A(fanout_net_42 ), .B1(_03415_ ), .B2(_03418_ ), .ZN(_01195_ ) );
NAND2_X1 _17416_ ( .A1(_03330_ ), .A2(_03174_ ), .ZN(_03419_ ) );
OAI21_X1 _17417_ ( .A(\u_lsu.pmem[3617] ), .B1(_03205_ ), .B2(_10532_ ), .ZN(_03420_ ) );
AOI21_X1 _17418_ ( .A(fanout_net_42 ), .B1(_03419_ ), .B2(_03420_ ), .ZN(_01196_ ) );
NAND4_X1 _17419_ ( .A1(_10402_ ), .A2(_03397_ ), .A3(_03407_ ), .A4(_03412_ ), .ZN(_03421_ ) );
OAI21_X1 _17420_ ( .A(\u_lsu.pmem[4774] ), .B1(_03405_ ), .B2(_03416_ ), .ZN(_03422_ ) );
AOI21_X1 _17421_ ( .A(fanout_net_42 ), .B1(_03421_ ), .B2(_03422_ ), .ZN(_01197_ ) );
NAND4_X1 _17422_ ( .A1(_10405_ ), .A2(_03397_ ), .A3(_03407_ ), .A4(_03412_ ), .ZN(_03423_ ) );
OAI21_X1 _17423_ ( .A(\u_lsu.pmem[4773] ), .B1(_03405_ ), .B2(_03416_ ), .ZN(_03424_ ) );
AOI21_X1 _17424_ ( .A(fanout_net_42 ), .B1(_03423_ ), .B2(_03424_ ), .ZN(_01198_ ) );
BUF_X4 _17425_ ( .A(_03396_ ), .Z(_03425_ ) );
NAND4_X1 _17426_ ( .A1(_10408_ ), .A2(_03425_ ), .A3(_03407_ ), .A4(_03412_ ), .ZN(_03426_ ) );
OAI21_X1 _17427_ ( .A(\u_lsu.pmem[4772] ), .B1(_03405_ ), .B2(_03416_ ), .ZN(_03427_ ) );
AOI21_X1 _17428_ ( .A(fanout_net_42 ), .B1(_03426_ ), .B2(_03427_ ), .ZN(_01199_ ) );
NAND4_X1 _17429_ ( .A1(_10411_ ), .A2(_03425_ ), .A3(_03407_ ), .A4(_03412_ ), .ZN(_03428_ ) );
OAI21_X1 _17430_ ( .A(\u_lsu.pmem[4771] ), .B1(_03405_ ), .B2(_03416_ ), .ZN(_03429_ ) );
AOI21_X1 _17431_ ( .A(fanout_net_42 ), .B1(_03428_ ), .B2(_03429_ ), .ZN(_01200_ ) );
NAND4_X1 _17432_ ( .A1(_10414_ ), .A2(_03425_ ), .A3(_03407_ ), .A4(_03412_ ), .ZN(_03430_ ) );
OAI21_X1 _17433_ ( .A(\u_lsu.pmem[4770] ), .B1(_03405_ ), .B2(_03416_ ), .ZN(_03431_ ) );
AOI21_X1 _17434_ ( .A(fanout_net_42 ), .B1(_03430_ ), .B2(_03431_ ), .ZN(_01201_ ) );
NAND4_X1 _17435_ ( .A1(_10417_ ), .A2(_03425_ ), .A3(_03407_ ), .A4(_03412_ ), .ZN(_03432_ ) );
BUF_X4 _17436_ ( .A(_09443_ ), .Z(_03433_ ) );
OAI21_X1 _17437_ ( .A(\u_lsu.pmem[4769] ), .B1(_03433_ ), .B2(_03416_ ), .ZN(_03434_ ) );
AOI21_X1 _17438_ ( .A(fanout_net_42 ), .B1(_03432_ ), .B2(_03434_ ), .ZN(_01202_ ) );
OAI21_X1 _17439_ ( .A(\u_lsu.pmem[4768] ), .B1(_03367_ ), .B2(_03417_ ), .ZN(_03435_ ) );
BUF_X4 _17440_ ( .A(_02484_ ), .Z(_03436_ ) );
NAND4_X1 _17441_ ( .A1(_02720_ ), .A2(_03242_ ), .A3(_03436_ ), .A4(_11292_ ), .ZN(_03437_ ) );
AOI21_X1 _17442_ ( .A(fanout_net_42 ), .B1(_03435_ ), .B2(_03437_ ), .ZN(_01203_ ) );
NAND3_X1 _17443_ ( .A1(_10423_ ), .A2(_02484_ ), .A3(_09842_ ), .ZN(_03438_ ) );
BUF_X4 _17444_ ( .A(_03438_ ), .Z(_03439_ ) );
BUF_X4 _17445_ ( .A(_10901_ ), .Z(_03440_ ) );
OAI21_X1 _17446_ ( .A(\u_lsu.pmem[4743] ), .B1(_03439_ ), .B2(_03440_ ), .ZN(_03441_ ) );
NAND4_X1 _17447_ ( .A1(_10436_ ), .A2(_03361_ ), .A3(_03371_ ), .A4(_03267_ ), .ZN(_03442_ ) );
AOI21_X1 _17448_ ( .A(fanout_net_42 ), .B1(_03441_ ), .B2(_03442_ ), .ZN(_01204_ ) );
BUF_X4 _17449_ ( .A(_03326_ ), .Z(_03443_ ) );
NAND4_X1 _17450_ ( .A1(_11321_ ), .A2(_09658_ ), .A3(_03443_ ), .A4(_03412_ ), .ZN(_03444_ ) );
OAI21_X1 _17451_ ( .A(\u_lsu.pmem[4742] ), .B1(_03439_ ), .B2(_02694_ ), .ZN(_03445_ ) );
AOI21_X1 _17452_ ( .A(fanout_net_42 ), .B1(_03444_ ), .B2(_03445_ ), .ZN(_01205_ ) );
NAND4_X1 _17453_ ( .A1(_11321_ ), .A2(_09713_ ), .A3(_02500_ ), .A4(_03412_ ), .ZN(_03446_ ) );
OAI21_X1 _17454_ ( .A(\u_lsu.pmem[4741] ), .B1(_03439_ ), .B2(_02694_ ), .ZN(_03447_ ) );
AOI21_X1 _17455_ ( .A(fanout_net_42 ), .B1(_03446_ ), .B2(_03447_ ), .ZN(_01206_ ) );
NAND4_X1 _17456_ ( .A1(_10556_ ), .A2(_03133_ ), .A3(_03299_ ), .A4(_03233_ ), .ZN(_03448_ ) );
OAI21_X1 _17457_ ( .A(\u_lsu.pmem[3616] ), .B1(_03205_ ), .B2(_10532_ ), .ZN(_03449_ ) );
AOI21_X1 _17458_ ( .A(fanout_net_42 ), .B1(_03448_ ), .B2(_03449_ ), .ZN(_01207_ ) );
BUF_X4 _17459_ ( .A(_03129_ ), .Z(_03450_ ) );
NAND4_X1 _17460_ ( .A1(_11321_ ), .A2(_09514_ ), .A3(_03443_ ), .A4(_03450_ ), .ZN(_03451_ ) );
OAI21_X1 _17461_ ( .A(\u_lsu.pmem[4740] ), .B1(_03439_ ), .B2(_02694_ ), .ZN(_03452_ ) );
AOI21_X1 _17462_ ( .A(fanout_net_42 ), .B1(_03451_ ), .B2(_03452_ ), .ZN(_01208_ ) );
NAND4_X1 _17463_ ( .A1(_11321_ ), .A2(_10456_ ), .A3(_02500_ ), .A4(_03450_ ), .ZN(_03453_ ) );
OAI21_X1 _17464_ ( .A(\u_lsu.pmem[4739] ), .B1(_03439_ ), .B2(_02694_ ), .ZN(_03454_ ) );
AOI21_X1 _17465_ ( .A(fanout_net_42 ), .B1(_03453_ ), .B2(_03454_ ), .ZN(_01209_ ) );
OAI21_X1 _17466_ ( .A(\u_lsu.pmem[4738] ), .B1(_03439_ ), .B2(_03440_ ), .ZN(_03455_ ) );
NAND4_X1 _17467_ ( .A1(_10460_ ), .A2(_03361_ ), .A3(_03371_ ), .A4(_03267_ ), .ZN(_03456_ ) );
AOI21_X1 _17468_ ( .A(fanout_net_42 ), .B1(_03455_ ), .B2(_03456_ ), .ZN(_01210_ ) );
BUF_X4 _17469_ ( .A(_11320_ ), .Z(_03457_ ) );
NAND4_X1 _17470_ ( .A1(_03457_ ), .A2(_09544_ ), .A3(_02500_ ), .A4(_03450_ ), .ZN(_03458_ ) );
OAI21_X1 _17471_ ( .A(\u_lsu.pmem[4737] ), .B1(_03439_ ), .B2(_09516_ ), .ZN(_03459_ ) );
AOI21_X1 _17472_ ( .A(fanout_net_42 ), .B1(_03458_ ), .B2(_03459_ ), .ZN(_01211_ ) );
NAND4_X1 _17473_ ( .A1(_03457_ ), .A2(_10467_ ), .A3(_02500_ ), .A4(_03450_ ), .ZN(_03460_ ) );
OAI21_X1 _17474_ ( .A(\u_lsu.pmem[4736] ), .B1(_03439_ ), .B2(_09516_ ), .ZN(_03461_ ) );
AOI21_X1 _17475_ ( .A(fanout_net_43 ), .B1(_03460_ ), .B2(_03461_ ), .ZN(_01212_ ) );
AND2_X2 _17476_ ( .A1(_11341_ ), .A2(_02409_ ), .ZN(_03462_ ) );
INV_X1 _17477_ ( .A(_03462_ ), .ZN(_03463_ ) );
BUF_X4 _17478_ ( .A(_03463_ ), .Z(_03464_ ) );
OAI21_X1 _17479_ ( .A(\u_lsu.pmem[4711] ), .B1(_03464_ ), .B2(_03440_ ), .ZN(_03465_ ) );
BUF_X4 _17480_ ( .A(_03462_ ), .Z(_03466_ ) );
NAND3_X1 _17481_ ( .A1(_11000_ ), .A2(_03466_ ), .A3(_11426_ ), .ZN(_03467_ ) );
AOI21_X1 _17482_ ( .A(fanout_net_43 ), .B1(_03465_ ), .B2(_03467_ ), .ZN(_01213_ ) );
OAI21_X1 _17483_ ( .A(\u_lsu.pmem[4710] ), .B1(_03464_ ), .B2(_03440_ ), .ZN(_03468_ ) );
NAND3_X1 _17484_ ( .A1(_10719_ ), .A2(_03466_ ), .A3(_11426_ ), .ZN(_03469_ ) );
AOI21_X1 _17485_ ( .A(fanout_net_43 ), .B1(_03468_ ), .B2(_03469_ ), .ZN(_01214_ ) );
OAI21_X1 _17486_ ( .A(\u_lsu.pmem[4709] ), .B1(_03464_ ), .B2(_03440_ ), .ZN(_03470_ ) );
NAND3_X1 _17487_ ( .A1(_10728_ ), .A2(_03466_ ), .A3(_11426_ ), .ZN(_03471_ ) );
AOI21_X1 _17488_ ( .A(fanout_net_43 ), .B1(_03470_ ), .B2(_03471_ ), .ZN(_01215_ ) );
OAI21_X1 _17489_ ( .A(\u_lsu.pmem[4708] ), .B1(_03464_ ), .B2(_03440_ ), .ZN(_03472_ ) );
BUF_X4 _17490_ ( .A(_09472_ ), .Z(_03473_ ) );
NAND3_X1 _17491_ ( .A1(_11152_ ), .A2(_03466_ ), .A3(_03473_ ), .ZN(_03474_ ) );
AOI21_X1 _17492_ ( .A(fanout_net_43 ), .B1(_03472_ ), .B2(_03474_ ), .ZN(_01216_ ) );
OAI21_X1 _17493_ ( .A(\u_lsu.pmem[4707] ), .B1(_03464_ ), .B2(_03440_ ), .ZN(_03475_ ) );
NAND3_X1 _17494_ ( .A1(_10733_ ), .A2(_03466_ ), .A3(_03473_ ), .ZN(_03476_ ) );
AOI21_X1 _17495_ ( .A(fanout_net_43 ), .B1(_03475_ ), .B2(_03476_ ), .ZN(_01217_ ) );
BUF_X2 _17496_ ( .A(_10041_ ), .Z(\alu_result_out[9] ) );
OAI21_X1 _17497_ ( .A(\u_lsu.pmem[3591] ), .B1(_10564_ ), .B2(\alu_result_out[9] ), .ZN(_03477_ ) );
BUF_X4 _17498_ ( .A(_08582_ ), .Z(_03478_ ) );
NAND4_X1 _17499_ ( .A1(_10566_ ), .A2(_03478_ ), .A3(_09496_ ), .A4(_09606_ ), .ZN(_03479_ ) );
AOI21_X1 _17500_ ( .A(fanout_net_43 ), .B1(_03477_ ), .B2(_03479_ ), .ZN(_01218_ ) );
OAI21_X1 _17501_ ( .A(\u_lsu.pmem[4706] ), .B1(_03464_ ), .B2(_03440_ ), .ZN(_03480_ ) );
NAND3_X1 _17502_ ( .A1(_09612_ ), .A2(_03466_ ), .A3(_03473_ ), .ZN(_03481_ ) );
AOI21_X1 _17503_ ( .A(fanout_net_43 ), .B1(_03480_ ), .B2(_03481_ ), .ZN(_01219_ ) );
OAI21_X1 _17504_ ( .A(\u_lsu.pmem[4705] ), .B1(_03464_ ), .B2(_03440_ ), .ZN(_03482_ ) );
NAND3_X1 _17505_ ( .A1(_10738_ ), .A2(_03466_ ), .A3(_03473_ ), .ZN(_03483_ ) );
AOI21_X1 _17506_ ( .A(fanout_net_43 ), .B1(_03482_ ), .B2(_03483_ ), .ZN(_01220_ ) );
OAI21_X1 _17507_ ( .A(\u_lsu.pmem[4704] ), .B1(_03464_ ), .B2(_03440_ ), .ZN(_03484_ ) );
NAND3_X1 _17508_ ( .A1(_10741_ ), .A2(_03466_ ), .A3(_03473_ ), .ZN(_03485_ ) );
AOI21_X1 _17509_ ( .A(fanout_net_43 ), .B1(_03484_ ), .B2(_03485_ ), .ZN(_01221_ ) );
AND2_X1 _17510_ ( .A1(_11369_ ), .A2(_09454_ ), .ZN(_03486_ ) );
INV_X1 _17511_ ( .A(_03486_ ), .ZN(_03487_ ) );
BUF_X4 _17512_ ( .A(_03487_ ), .Z(_03488_ ) );
BUF_X4 _17513_ ( .A(_10901_ ), .Z(_03489_ ) );
OAI21_X1 _17514_ ( .A(\u_lsu.pmem[4679] ), .B1(_03488_ ), .B2(_03489_ ), .ZN(_03490_ ) );
NAND4_X1 _17515_ ( .A1(_09742_ ), .A2(_03242_ ), .A3(_03371_ ), .A4(_11378_ ), .ZN(_03491_ ) );
AOI21_X1 _17516_ ( .A(fanout_net_43 ), .B1(_03490_ ), .B2(_03491_ ), .ZN(_01222_ ) );
OAI21_X1 _17517_ ( .A(\u_lsu.pmem[4678] ), .B1(_03488_ ), .B2(_03489_ ), .ZN(_03492_ ) );
NAND4_X1 _17518_ ( .A1(_11347_ ), .A2(_03242_ ), .A3(_03371_ ), .A4(_11378_ ), .ZN(_03493_ ) );
AOI21_X1 _17519_ ( .A(fanout_net_43 ), .B1(_03492_ ), .B2(_03493_ ), .ZN(_01223_ ) );
OAI21_X1 _17520_ ( .A(\u_lsu.pmem[4677] ), .B1(_03488_ ), .B2(_03489_ ), .ZN(_03494_ ) );
NAND4_X1 _17521_ ( .A1(_11351_ ), .A2(_03242_ ), .A3(_03371_ ), .A4(_11378_ ), .ZN(_03495_ ) );
AOI21_X1 _17522_ ( .A(fanout_net_43 ), .B1(_03494_ ), .B2(_03495_ ), .ZN(_01224_ ) );
OAI21_X1 _17523_ ( .A(\u_lsu.pmem[4676] ), .B1(_03488_ ), .B2(_03489_ ), .ZN(_03496_ ) );
NAND4_X1 _17524_ ( .A1(_02327_ ), .A2(_03242_ ), .A3(_03371_ ), .A4(_11378_ ), .ZN(_03497_ ) );
AOI21_X1 _17525_ ( .A(fanout_net_43 ), .B1(_03496_ ), .B2(_03497_ ), .ZN(_01225_ ) );
OAI21_X1 _17526_ ( .A(\u_lsu.pmem[4675] ), .B1(_03488_ ), .B2(_03489_ ), .ZN(_03498_ ) );
BUF_X4 _17527_ ( .A(_11369_ ), .Z(_03499_ ) );
NAND4_X1 _17528_ ( .A1(_03091_ ), .A2(_03242_ ), .A3(_03371_ ), .A4(_03499_ ), .ZN(_03500_ ) );
AOI21_X1 _17529_ ( .A(fanout_net_43 ), .B1(_03498_ ), .B2(_03500_ ), .ZN(_01226_ ) );
OAI21_X1 _17530_ ( .A(\u_lsu.pmem[4674] ), .B1(_03488_ ), .B2(_03489_ ), .ZN(_03501_ ) );
NAND4_X1 _17531_ ( .A1(_02379_ ), .A2(_03242_ ), .A3(_03371_ ), .A4(_03499_ ), .ZN(_03502_ ) );
AOI21_X1 _17532_ ( .A(fanout_net_43 ), .B1(_03501_ ), .B2(_03502_ ), .ZN(_01227_ ) );
OAI21_X1 _17533_ ( .A(\u_lsu.pmem[4673] ), .B1(_03488_ ), .B2(_03489_ ), .ZN(_03503_ ) );
BUF_X4 _17534_ ( .A(_09950_ ), .Z(_03504_ ) );
BUF_X4 _17535_ ( .A(_02881_ ), .Z(_03505_ ) );
NAND4_X1 _17536_ ( .A1(_03143_ ), .A2(_03504_ ), .A3(_03505_ ), .A4(_03499_ ), .ZN(_03506_ ) );
AOI21_X1 _17537_ ( .A(fanout_net_43 ), .B1(_03503_ ), .B2(_03506_ ), .ZN(_01228_ ) );
OAI21_X1 _17538_ ( .A(\u_lsu.pmem[3590] ), .B1(_10564_ ), .B2(\alu_result_out[9] ), .ZN(_03507_ ) );
NAND4_X1 _17539_ ( .A1(_10566_ ), .A2(_03056_ ), .A3(_09496_ ), .A4(_09606_ ), .ZN(_03508_ ) );
AOI21_X1 _17540_ ( .A(fanout_net_43 ), .B1(_03507_ ), .B2(_03508_ ), .ZN(_01229_ ) );
OAI21_X1 _17541_ ( .A(\u_lsu.pmem[4672] ), .B1(_03488_ ), .B2(_03489_ ), .ZN(_03509_ ) );
NAND4_X1 _17542_ ( .A1(_02720_ ), .A2(_03504_ ), .A3(_03505_ ), .A4(_03499_ ), .ZN(_03510_ ) );
AOI21_X1 _17543_ ( .A(fanout_net_43 ), .B1(_03509_ ), .B2(_03510_ ), .ZN(_01230_ ) );
NAND4_X1 _17544_ ( .A1(_10527_ ), .A2(_03425_ ), .A3(_03443_ ), .A4(_03450_ ), .ZN(_03511_ ) );
AND3_X2 _17545_ ( .A1(_09538_ ), .A2(_02409_ ), .A3(_10530_ ), .ZN(_03512_ ) );
INV_X1 _17546_ ( .A(_03512_ ), .ZN(_03513_ ) );
OAI21_X1 _17547_ ( .A(\u_lsu.pmem[4647] ), .B1(_03433_ ), .B2(_03513_ ), .ZN(_03514_ ) );
AOI21_X1 _17548_ ( .A(fanout_net_43 ), .B1(_03511_ ), .B2(_03514_ ), .ZN(_01231_ ) );
NAND4_X1 _17549_ ( .A1(_10535_ ), .A2(_03425_ ), .A3(_03443_ ), .A4(_03450_ ), .ZN(_03515_ ) );
OAI21_X1 _17550_ ( .A(\u_lsu.pmem[4646] ), .B1(_03433_ ), .B2(_03513_ ), .ZN(_03516_ ) );
AOI21_X1 _17551_ ( .A(fanout_net_43 ), .B1(_03515_ ), .B2(_03516_ ), .ZN(_01232_ ) );
NAND4_X1 _17552_ ( .A1(_10538_ ), .A2(_03425_ ), .A3(_03443_ ), .A4(_03450_ ), .ZN(_03517_ ) );
OAI21_X1 _17553_ ( .A(\u_lsu.pmem[4645] ), .B1(_03433_ ), .B2(_03513_ ), .ZN(_03518_ ) );
AOI21_X1 _17554_ ( .A(fanout_net_43 ), .B1(_03517_ ), .B2(_03518_ ), .ZN(_01233_ ) );
BUF_X4 _17555_ ( .A(_03513_ ), .Z(_03519_ ) );
OAI21_X1 _17556_ ( .A(\u_lsu.pmem[4644] ), .B1(_03367_ ), .B2(_03519_ ), .ZN(_03520_ ) );
NAND3_X1 _17557_ ( .A1(_11152_ ), .A2(_03306_ ), .A3(_03512_ ), .ZN(_03521_ ) );
AOI21_X1 _17558_ ( .A(fanout_net_43 ), .B1(_03520_ ), .B2(_03521_ ), .ZN(_01234_ ) );
OAI21_X1 _17559_ ( .A(\u_lsu.pmem[4643] ), .B1(_03367_ ), .B2(_03519_ ), .ZN(_03522_ ) );
NAND3_X1 _17560_ ( .A1(_10733_ ), .A2(_11214_ ), .A3(_03512_ ), .ZN(_03523_ ) );
AOI21_X1 _17561_ ( .A(fanout_net_43 ), .B1(_03522_ ), .B2(_03523_ ), .ZN(_01235_ ) );
OAI21_X1 _17562_ ( .A(\u_lsu.pmem[4642] ), .B1(_03367_ ), .B2(_03513_ ), .ZN(_03524_ ) );
NAND3_X1 _17563_ ( .A1(_09612_ ), .A2(_03512_ ), .A3(_03473_ ), .ZN(_03525_ ) );
AOI21_X1 _17564_ ( .A(fanout_net_43 ), .B1(_03524_ ), .B2(_03525_ ), .ZN(_01236_ ) );
OAI21_X1 _17565_ ( .A(\u_lsu.pmem[4641] ), .B1(_03367_ ), .B2(_03513_ ), .ZN(_03526_ ) );
NAND3_X1 _17566_ ( .A1(_10738_ ), .A2(_11214_ ), .A3(_03512_ ), .ZN(_03527_ ) );
AOI21_X1 _17567_ ( .A(fanout_net_43 ), .B1(_03526_ ), .B2(_03527_ ), .ZN(_01237_ ) );
NAND4_X1 _17568_ ( .A1(_10556_ ), .A2(_03425_ ), .A3(_03443_ ), .A4(_03450_ ), .ZN(_03528_ ) );
OAI21_X1 _17569_ ( .A(\u_lsu.pmem[4640] ), .B1(_03433_ ), .B2(_03513_ ), .ZN(_03529_ ) );
AOI21_X1 _17570_ ( .A(fanout_net_43 ), .B1(_03528_ ), .B2(_03529_ ), .ZN(_01238_ ) );
AND3_X1 _17571_ ( .A1(_09453_ ), .A2(_10560_ ), .A3(_09538_ ), .ZN(_03530_ ) );
INV_X1 _17572_ ( .A(_03530_ ), .ZN(_03531_ ) );
BUF_X4 _17573_ ( .A(_03531_ ), .Z(_03532_ ) );
OAI21_X1 _17574_ ( .A(\u_lsu.pmem[4615] ), .B1(_03532_ ), .B2(_03489_ ), .ZN(_03533_ ) );
BUF_X4 _17575_ ( .A(_03530_ ), .Z(_03534_ ) );
NAND3_X1 _17576_ ( .A1(_03534_ ), .A2(_11423_ ), .A3(_03473_ ), .ZN(_03535_ ) );
AOI21_X1 _17577_ ( .A(fanout_net_43 ), .B1(_03533_ ), .B2(_03535_ ), .ZN(_01239_ ) );
OAI21_X1 _17578_ ( .A(\u_lsu.pmem[3589] ), .B1(_10564_ ), .B2(\alu_result_out[9] ), .ZN(_03536_ ) );
NAND4_X1 _17579_ ( .A1(_10566_ ), .A2(_03059_ ), .A3(_09496_ ), .A4(_09606_ ), .ZN(_03537_ ) );
AOI21_X1 _17580_ ( .A(fanout_net_43 ), .B1(_03536_ ), .B2(_03537_ ), .ZN(_01240_ ) );
OAI21_X1 _17581_ ( .A(\u_lsu.pmem[4614] ), .B1(_03532_ ), .B2(_03489_ ), .ZN(_03538_ ) );
NAND3_X1 _17582_ ( .A1(_03534_ ), .A2(_10444_ ), .A3(_03473_ ), .ZN(_03539_ ) );
AOI21_X1 _17583_ ( .A(fanout_net_43 ), .B1(_03538_ ), .B2(_03539_ ), .ZN(_01241_ ) );
BUF_X4 _17584_ ( .A(_09675_ ), .Z(_03540_ ) );
OAI21_X1 _17585_ ( .A(\u_lsu.pmem[4613] ), .B1(_03532_ ), .B2(_03540_ ), .ZN(_03541_ ) );
NAND3_X1 _17586_ ( .A1(_03534_ ), .A2(_10448_ ), .A3(_03473_ ), .ZN(_03542_ ) );
AOI21_X1 _17587_ ( .A(fanout_net_44 ), .B1(_03541_ ), .B2(_03542_ ), .ZN(_01242_ ) );
OAI21_X1 _17588_ ( .A(\u_lsu.pmem[4612] ), .B1(_03532_ ), .B2(_03540_ ), .ZN(_03543_ ) );
NAND3_X1 _17589_ ( .A1(_03534_ ), .A2(_10453_ ), .A3(_03473_ ), .ZN(_03544_ ) );
AOI21_X1 _17590_ ( .A(fanout_net_44 ), .B1(_03543_ ), .B2(_03544_ ), .ZN(_01243_ ) );
NAND4_X1 _17591_ ( .A1(_10575_ ), .A2(_03425_ ), .A3(_03443_ ), .A4(_03450_ ), .ZN(_03545_ ) );
OAI21_X1 _17592_ ( .A(\u_lsu.pmem[4611] ), .B1(_03531_ ), .B2(_09516_ ), .ZN(_03546_ ) );
AOI21_X1 _17593_ ( .A(fanout_net_44 ), .B1(_03545_ ), .B2(_03546_ ), .ZN(_01244_ ) );
NAND4_X1 _17594_ ( .A1(_10584_ ), .A2(_09806_ ), .A3(_03443_ ), .A4(_03450_ ), .ZN(_03547_ ) );
OAI21_X1 _17595_ ( .A(\u_lsu.pmem[4610] ), .B1(_03531_ ), .B2(_09516_ ), .ZN(_03548_ ) );
AOI21_X1 _17596_ ( .A(fanout_net_44 ), .B1(_03547_ ), .B2(_03548_ ), .ZN(_01245_ ) );
OAI21_X1 _17597_ ( .A(\u_lsu.pmem[4609] ), .B1(_03532_ ), .B2(_03540_ ), .ZN(_03549_ ) );
BUF_X4 _17598_ ( .A(_09472_ ), .Z(_03550_ ) );
NAND3_X1 _17599_ ( .A1(_03534_ ), .A2(_10463_ ), .A3(_03550_ ), .ZN(_03551_ ) );
AOI21_X1 _17600_ ( .A(fanout_net_44 ), .B1(_03549_ ), .B2(_03551_ ), .ZN(_01246_ ) );
BUF_X4 _17601_ ( .A(_03129_ ), .Z(_03552_ ) );
NAND4_X1 _17602_ ( .A1(_10591_ ), .A2(_03425_ ), .A3(_03443_ ), .A4(_03552_ ), .ZN(_03553_ ) );
OAI21_X1 _17603_ ( .A(\u_lsu.pmem[4608] ), .B1(_03531_ ), .B2(_09516_ ), .ZN(_03554_ ) );
AOI21_X1 _17604_ ( .A(fanout_net_44 ), .B1(_03553_ ), .B2(_03554_ ), .ZN(_01247_ ) );
NAND2_X1 _17605_ ( .A1(_02980_ ), .A2(_11442_ ), .ZN(_03555_ ) );
BUF_X4 _17606_ ( .A(_03555_ ), .Z(_03556_ ) );
OAI21_X1 _17607_ ( .A(\u_lsu.pmem[4583] ), .B1(_03367_ ), .B2(_03556_ ), .ZN(_03557_ ) );
NAND4_X1 _17608_ ( .A1(_09742_ ), .A2(_03504_ ), .A3(_03505_ ), .A4(_11442_ ), .ZN(_03558_ ) );
AOI21_X1 _17609_ ( .A(fanout_net_44 ), .B1(_03557_ ), .B2(_03558_ ), .ZN(_01248_ ) );
BUF_X4 _17610_ ( .A(_03396_ ), .Z(_03559_ ) );
NAND4_X1 _17611_ ( .A1(_10603_ ), .A2(_03559_ ), .A3(_03443_ ), .A4(_03552_ ), .ZN(_03560_ ) );
OAI21_X1 _17612_ ( .A(\u_lsu.pmem[4582] ), .B1(_03433_ ), .B2(_03556_ ), .ZN(_03561_ ) );
AOI21_X1 _17613_ ( .A(fanout_net_44 ), .B1(_03560_ ), .B2(_03561_ ), .ZN(_01249_ ) );
BUF_X4 _17614_ ( .A(_03326_ ), .Z(_03562_ ) );
NAND4_X1 _17615_ ( .A1(_10608_ ), .A2(_03559_ ), .A3(_03562_ ), .A4(_03552_ ), .ZN(_03563_ ) );
OAI21_X1 _17616_ ( .A(\u_lsu.pmem[4581] ), .B1(_03433_ ), .B2(_03555_ ), .ZN(_03564_ ) );
AOI21_X1 _17617_ ( .A(fanout_net_44 ), .B1(_03563_ ), .B2(_03564_ ), .ZN(_01250_ ) );
OAI21_X1 _17618_ ( .A(\u_lsu.pmem[4386] ), .B1(_09441_ ), .B2(_03540_ ), .ZN(_03565_ ) );
NAND4_X1 _17619_ ( .A1(_09938_ ), .A2(_03504_ ), .A3(_09131_ ), .A4(_09456_ ), .ZN(_03566_ ) );
AOI21_X1 _17620_ ( .A(fanout_net_44 ), .B1(_03565_ ), .B2(_03566_ ), .ZN(_01251_ ) );
NAND4_X1 _17621_ ( .A1(_09791_ ), .A2(_03559_ ), .A3(_03562_ ), .A4(_03552_ ), .ZN(_03567_ ) );
OAI21_X1 _17622_ ( .A(\u_lsu.pmem[4320] ), .B1(_03433_ ), .B2(_09751_ ), .ZN(_03568_ ) );
AOI21_X1 _17623_ ( .A(fanout_net_44 ), .B1(_03567_ ), .B2(_03568_ ), .ZN(_01252_ ) );
OAI21_X1 _17624_ ( .A(\u_lsu.pmem[3588] ), .B1(_10564_ ), .B2(\alu_result_out[9] ), .ZN(_03569_ ) );
NAND4_X1 _17625_ ( .A1(_10566_ ), .A2(_03064_ ), .A3(_09496_ ), .A4(_09606_ ), .ZN(_03570_ ) );
AOI21_X1 _17626_ ( .A(fanout_net_44 ), .B1(_03569_ ), .B2(_03570_ ), .ZN(_01253_ ) );
NAND4_X1 _17627_ ( .A1(_10611_ ), .A2(_03559_ ), .A3(_03562_ ), .A4(_03552_ ), .ZN(_03571_ ) );
OAI21_X1 _17628_ ( .A(\u_lsu.pmem[4580] ), .B1(_03433_ ), .B2(_03555_ ), .ZN(_03572_ ) );
AOI21_X1 _17629_ ( .A(fanout_net_44 ), .B1(_03571_ ), .B2(_03572_ ), .ZN(_01254_ ) );
NAND4_X1 _17630_ ( .A1(_10614_ ), .A2(_03559_ ), .A3(_03562_ ), .A4(_03552_ ), .ZN(_03573_ ) );
OAI21_X1 _17631_ ( .A(\u_lsu.pmem[4579] ), .B1(_03433_ ), .B2(_03555_ ), .ZN(_03574_ ) );
AOI21_X1 _17632_ ( .A(fanout_net_44 ), .B1(_03573_ ), .B2(_03574_ ), .ZN(_01255_ ) );
NAND4_X1 _17633_ ( .A1(_10617_ ), .A2(_03559_ ), .A3(_03562_ ), .A4(_03552_ ), .ZN(_03575_ ) );
BUF_X4 _17634_ ( .A(_09443_ ), .Z(_03576_ ) );
OAI21_X1 _17635_ ( .A(\u_lsu.pmem[4578] ), .B1(_03576_ ), .B2(_03555_ ), .ZN(_03577_ ) );
AOI21_X1 _17636_ ( .A(fanout_net_44 ), .B1(_03575_ ), .B2(_03577_ ), .ZN(_01256_ ) );
NAND4_X1 _17637_ ( .A1(_10621_ ), .A2(_03559_ ), .A3(_03562_ ), .A4(_03552_ ), .ZN(_03578_ ) );
OAI21_X1 _17638_ ( .A(\u_lsu.pmem[4577] ), .B1(_03576_ ), .B2(_03555_ ), .ZN(_03579_ ) );
AOI21_X1 _17639_ ( .A(fanout_net_44 ), .B1(_03578_ ), .B2(_03579_ ), .ZN(_01257_ ) );
NAND4_X1 _17640_ ( .A1(_10624_ ), .A2(_03559_ ), .A3(_03562_ ), .A4(_03552_ ), .ZN(_03580_ ) );
OAI21_X1 _17641_ ( .A(\u_lsu.pmem[4576] ), .B1(_03576_ ), .B2(_03555_ ), .ZN(_03581_ ) );
AOI21_X1 _17642_ ( .A(fanout_net_44 ), .B1(_03580_ ), .B2(_03581_ ), .ZN(_01258_ ) );
NAND2_X1 _17643_ ( .A1(_02980_ ), .A2(_11469_ ), .ZN(_03582_ ) );
BUF_X4 _17644_ ( .A(_03582_ ), .Z(_03583_ ) );
OAI21_X1 _17645_ ( .A(\u_lsu.pmem[4551] ), .B1(_03367_ ), .B2(_03583_ ), .ZN(_03584_ ) );
NAND4_X1 _17646_ ( .A1(_09742_ ), .A2(_03504_ ), .A3(_03505_ ), .A4(_11469_ ), .ZN(_03585_ ) );
AOI21_X1 _17647_ ( .A(fanout_net_44 ), .B1(_03584_ ), .B2(_03585_ ), .ZN(_01259_ ) );
NAND4_X1 _17648_ ( .A1(_10632_ ), .A2(_03559_ ), .A3(_03562_ ), .A4(_03552_ ), .ZN(_03586_ ) );
OAI21_X1 _17649_ ( .A(\u_lsu.pmem[4550] ), .B1(_03576_ ), .B2(_03583_ ), .ZN(_03587_ ) );
AOI21_X1 _17650_ ( .A(fanout_net_44 ), .B1(_03586_ ), .B2(_03587_ ), .ZN(_01260_ ) );
BUF_X4 _17651_ ( .A(_03129_ ), .Z(_03588_ ) );
NAND4_X1 _17652_ ( .A1(_10635_ ), .A2(_03559_ ), .A3(_03562_ ), .A4(_03588_ ), .ZN(_03589_ ) );
OAI21_X1 _17653_ ( .A(\u_lsu.pmem[4549] ), .B1(_03576_ ), .B2(_03582_ ), .ZN(_03590_ ) );
AOI21_X1 _17654_ ( .A(fanout_net_44 ), .B1(_03589_ ), .B2(_03590_ ), .ZN(_01261_ ) );
BUF_X4 _17655_ ( .A(_03396_ ), .Z(_03591_ ) );
NAND4_X1 _17656_ ( .A1(_10641_ ), .A2(_03591_ ), .A3(_03562_ ), .A4(_03588_ ), .ZN(_03592_ ) );
OAI21_X1 _17657_ ( .A(\u_lsu.pmem[4548] ), .B1(_03576_ ), .B2(_03582_ ), .ZN(_03593_ ) );
AOI21_X1 _17658_ ( .A(fanout_net_44 ), .B1(_03592_ ), .B2(_03593_ ), .ZN(_01262_ ) );
BUF_X4 _17659_ ( .A(_03326_ ), .Z(_03594_ ) );
NAND4_X1 _17660_ ( .A1(_10645_ ), .A2(_03591_ ), .A3(_03594_ ), .A4(_03588_ ), .ZN(_03595_ ) );
OAI21_X1 _17661_ ( .A(\u_lsu.pmem[4547] ), .B1(_03576_ ), .B2(_03582_ ), .ZN(_03596_ ) );
AOI21_X1 _17662_ ( .A(fanout_net_44 ), .B1(_03595_ ), .B2(_03596_ ), .ZN(_01263_ ) );
NAND4_X1 _17663_ ( .A1(_10575_ ), .A2(_02976_ ), .A3(_03299_ ), .A4(_03233_ ), .ZN(_03597_ ) );
OAI21_X1 _17664_ ( .A(\u_lsu.pmem[3587] ), .B1(_10563_ ), .B2(_10910_ ), .ZN(_03598_ ) );
AOI21_X1 _17665_ ( .A(fanout_net_44 ), .B1(_03597_ ), .B2(_03598_ ), .ZN(_01264_ ) );
NAND4_X1 _17666_ ( .A1(_10649_ ), .A2(_03591_ ), .A3(_03594_ ), .A4(_03588_ ), .ZN(_03599_ ) );
OAI21_X1 _17667_ ( .A(\u_lsu.pmem[4546] ), .B1(_03576_ ), .B2(_03582_ ), .ZN(_03600_ ) );
AOI21_X1 _17668_ ( .A(fanout_net_44 ), .B1(_03599_ ), .B2(_03600_ ), .ZN(_01265_ ) );
NAND4_X1 _17669_ ( .A1(_10652_ ), .A2(_03591_ ), .A3(_03594_ ), .A4(_03588_ ), .ZN(_03601_ ) );
OAI21_X1 _17670_ ( .A(\u_lsu.pmem[4545] ), .B1(_03576_ ), .B2(_03582_ ), .ZN(_03602_ ) );
AOI21_X1 _17671_ ( .A(fanout_net_44 ), .B1(_03601_ ), .B2(_03602_ ), .ZN(_01266_ ) );
NAND4_X1 _17672_ ( .A1(_10655_ ), .A2(_03591_ ), .A3(_03594_ ), .A4(_03588_ ), .ZN(_03603_ ) );
OAI21_X1 _17673_ ( .A(\u_lsu.pmem[4544] ), .B1(_03576_ ), .B2(_03582_ ), .ZN(_03604_ ) );
AOI21_X1 _17674_ ( .A(fanout_net_44 ), .B1(_03603_ ), .B2(_03604_ ), .ZN(_01267_ ) );
NAND4_X1 _17675_ ( .A1(_10658_ ), .A2(_03591_ ), .A3(_03594_ ), .A4(_03588_ ), .ZN(_03605_ ) );
BUF_X4 _17676_ ( .A(_09443_ ), .Z(_03606_ ) );
NAND2_X1 _17677_ ( .A1(_11499_ ), .A2(_02980_ ), .ZN(_03607_ ) );
BUF_X4 _17678_ ( .A(_03607_ ), .Z(_03608_ ) );
OAI21_X1 _17679_ ( .A(\u_lsu.pmem[4519] ), .B1(_03606_ ), .B2(_03608_ ), .ZN(_03609_ ) );
AOI21_X1 _17680_ ( .A(fanout_net_44 ), .B1(_03605_ ), .B2(_03609_ ), .ZN(_01268_ ) );
NAND4_X1 _17681_ ( .A1(_10665_ ), .A2(_03591_ ), .A3(_03594_ ), .A4(_03588_ ), .ZN(_03610_ ) );
OAI21_X1 _17682_ ( .A(\u_lsu.pmem[4518] ), .B1(_03606_ ), .B2(_03607_ ), .ZN(_03611_ ) );
AOI21_X1 _17683_ ( .A(fanout_net_44 ), .B1(_03610_ ), .B2(_03611_ ), .ZN(_01269_ ) );
NAND4_X1 _17684_ ( .A1(_10668_ ), .A2(_03591_ ), .A3(_03594_ ), .A4(_03588_ ), .ZN(_03612_ ) );
OAI21_X1 _17685_ ( .A(\u_lsu.pmem[4517] ), .B1(_03606_ ), .B2(_03607_ ), .ZN(_03613_ ) );
AOI21_X1 _17686_ ( .A(fanout_net_44 ), .B1(_03612_ ), .B2(_03613_ ), .ZN(_01270_ ) );
NAND4_X1 _17687_ ( .A1(_10671_ ), .A2(_03591_ ), .A3(_03594_ ), .A4(_03588_ ), .ZN(_03614_ ) );
OAI21_X1 _17688_ ( .A(\u_lsu.pmem[4516] ), .B1(_03606_ ), .B2(_03607_ ), .ZN(_03615_ ) );
AOI21_X1 _17689_ ( .A(fanout_net_44 ), .B1(_03614_ ), .B2(_03615_ ), .ZN(_01271_ ) );
BUF_X4 _17690_ ( .A(_03129_ ), .Z(_03616_ ) );
NAND4_X1 _17691_ ( .A1(_10674_ ), .A2(_03591_ ), .A3(_03594_ ), .A4(_03616_ ), .ZN(_03617_ ) );
OAI21_X1 _17692_ ( .A(\u_lsu.pmem[4515] ), .B1(_03606_ ), .B2(_03607_ ), .ZN(_03618_ ) );
AOI21_X1 _17693_ ( .A(fanout_net_45 ), .B1(_03617_ ), .B2(_03618_ ), .ZN(_01272_ ) );
BUF_X4 _17694_ ( .A(_03396_ ), .Z(_03619_ ) );
NAND4_X1 _17695_ ( .A1(_10679_ ), .A2(_03619_ ), .A3(_03594_ ), .A4(_03616_ ), .ZN(_03620_ ) );
OAI21_X1 _17696_ ( .A(\u_lsu.pmem[4514] ), .B1(_03606_ ), .B2(_03607_ ), .ZN(_03621_ ) );
AOI21_X1 _17697_ ( .A(fanout_net_45 ), .B1(_03620_ ), .B2(_03621_ ), .ZN(_01273_ ) );
BUF_X4 _17698_ ( .A(_03326_ ), .Z(_03622_ ) );
NAND4_X1 _17699_ ( .A1(_10682_ ), .A2(_03619_ ), .A3(_03622_ ), .A4(_03616_ ), .ZN(_03623_ ) );
OAI21_X1 _17700_ ( .A(\u_lsu.pmem[4513] ), .B1(_03606_ ), .B2(_03607_ ), .ZN(_03624_ ) );
AOI21_X1 _17701_ ( .A(fanout_net_45 ), .B1(_03623_ ), .B2(_03624_ ), .ZN(_01274_ ) );
NAND4_X1 _17702_ ( .A1(_10584_ ), .A2(_10974_ ), .A3(\alu_result_out[8] ), .A4(_10585_ ), .ZN(_03625_ ) );
OAI21_X1 _17703_ ( .A(\u_lsu.pmem[3586] ), .B1(_10563_ ), .B2(_10910_ ), .ZN(_03626_ ) );
AOI21_X1 _17704_ ( .A(fanout_net_45 ), .B1(_03625_ ), .B2(_03626_ ), .ZN(_01275_ ) );
OAI21_X1 _17705_ ( .A(\u_lsu.pmem[4512] ), .B1(_03367_ ), .B2(_03608_ ), .ZN(_03627_ ) );
NAND4_X1 _17706_ ( .A1(_02720_ ), .A2(_03504_ ), .A3(_03505_ ), .A4(_11499_ ), .ZN(_03628_ ) );
AOI21_X1 _17707_ ( .A(fanout_net_45 ), .B1(_03627_ ), .B2(_03628_ ), .ZN(_01276_ ) );
OAI21_X1 _17708_ ( .A(\u_lsu.pmem[4487] ), .B1(_09509_ ), .B2(_03540_ ), .ZN(_03629_ ) );
NAND4_X1 _17709_ ( .A1(_11542_ ), .A2(_03478_ ), .A3(_03505_ ), .A4(_03267_ ), .ZN(_03630_ ) );
AOI21_X1 _17710_ ( .A(fanout_net_45 ), .B1(_03629_ ), .B2(_03630_ ), .ZN(_01277_ ) );
OAI21_X1 _17711_ ( .A(\u_lsu.pmem[4486] ), .B1(_09509_ ), .B2(_03540_ ), .ZN(_03631_ ) );
NAND4_X1 _17712_ ( .A1(_11542_ ), .A2(_03056_ ), .A3(_03505_ ), .A4(_03267_ ), .ZN(_03632_ ) );
AOI21_X1 _17713_ ( .A(fanout_net_45 ), .B1(_03631_ ), .B2(_03632_ ), .ZN(_01278_ ) );
OAI21_X1 _17714_ ( .A(\u_lsu.pmem[4485] ), .B1(_09509_ ), .B2(_03540_ ), .ZN(_03633_ ) );
NAND4_X1 _17715_ ( .A1(_11542_ ), .A2(_03059_ ), .A3(_03505_ ), .A4(_03267_ ), .ZN(_03634_ ) );
AOI21_X1 _17716_ ( .A(fanout_net_45 ), .B1(_03633_ ), .B2(_03634_ ), .ZN(_01279_ ) );
OAI21_X1 _17717_ ( .A(\u_lsu.pmem[4484] ), .B1(_09509_ ), .B2(_03540_ ), .ZN(_03635_ ) );
NAND4_X1 _17718_ ( .A1(_11542_ ), .A2(_03064_ ), .A3(_03505_ ), .A4(_03267_ ), .ZN(_03636_ ) );
AOI21_X1 _17719_ ( .A(fanout_net_45 ), .B1(_03635_ ), .B2(_03636_ ), .ZN(_01280_ ) );
OAI21_X1 _17720_ ( .A(\u_lsu.pmem[4483] ), .B1(_09509_ ), .B2(_03540_ ), .ZN(_03637_ ) );
NAND4_X1 _17721_ ( .A1(_11542_ ), .A2(_10915_ ), .A3(_03505_ ), .A4(_03267_ ), .ZN(_03638_ ) );
AOI21_X1 _17722_ ( .A(fanout_net_45 ), .B1(_03637_ ), .B2(_03638_ ), .ZN(_01281_ ) );
OAI21_X1 _17723_ ( .A(\u_lsu.pmem[4482] ), .B1(_09508_ ), .B2(_03540_ ), .ZN(_03639_ ) );
BUF_X4 _17724_ ( .A(_02881_ ), .Z(_03640_ ) );
NAND4_X1 _17725_ ( .A1(_09537_ ), .A2(_03361_ ), .A3(_03640_ ), .A4(_03267_ ), .ZN(_03641_ ) );
AOI21_X1 _17726_ ( .A(fanout_net_45 ), .B1(_03639_ ), .B2(_03641_ ), .ZN(_01282_ ) );
BUF_X4 _17727_ ( .A(_09675_ ), .Z(_03642_ ) );
OAI21_X1 _17728_ ( .A(\u_lsu.pmem[4481] ), .B1(_09508_ ), .B2(_03642_ ), .ZN(_03643_ ) );
NAND4_X1 _17729_ ( .A1(_11542_ ), .A2(_02308_ ), .A3(_03640_ ), .A4(_03267_ ), .ZN(_03644_ ) );
AOI21_X1 _17730_ ( .A(fanout_net_45 ), .B1(_03643_ ), .B2(_03644_ ), .ZN(_01283_ ) );
OAI21_X1 _17731_ ( .A(\u_lsu.pmem[4480] ), .B1(_09508_ ), .B2(_03642_ ), .ZN(_03645_ ) );
BUF_X4 _17732_ ( .A(_10904_ ), .Z(_03646_ ) );
NAND4_X1 _17733_ ( .A1(_11542_ ), .A2(_11131_ ), .A3(_03640_ ), .A4(_03646_ ), .ZN(_03647_ ) );
AOI21_X1 _17734_ ( .A(fanout_net_45 ), .B1(_03645_ ), .B2(_03647_ ), .ZN(_01284_ ) );
OAI21_X1 _17735_ ( .A(\u_lsu.pmem[4455] ), .B1(_09569_ ), .B2(_03642_ ), .ZN(_03648_ ) );
NAND3_X1 _17736_ ( .A1(_11000_ ), .A2(_09574_ ), .A3(_03550_ ), .ZN(_03649_ ) );
AOI21_X1 _17737_ ( .A(fanout_net_45 ), .B1(_03648_ ), .B2(_03649_ ), .ZN(_01285_ ) );
OAI21_X1 _17738_ ( .A(\u_lsu.pmem[3585] ), .B1(_10564_ ), .B2(\alu_result_out[9] ), .ZN(_03650_ ) );
NAND4_X1 _17739_ ( .A1(_10566_ ), .A2(_02308_ ), .A3(_09496_ ), .A4(_09606_ ), .ZN(_03651_ ) );
AOI21_X1 _17740_ ( .A(fanout_net_45 ), .B1(_03650_ ), .B2(_03651_ ), .ZN(_01286_ ) );
OAI21_X1 _17741_ ( .A(\u_lsu.pmem[4454] ), .B1(_09569_ ), .B2(_03642_ ), .ZN(_03652_ ) );
NAND3_X1 _17742_ ( .A1(_10719_ ), .A2(_09574_ ), .A3(_03550_ ), .ZN(_03653_ ) );
AOI21_X1 _17743_ ( .A(fanout_net_45 ), .B1(_03652_ ), .B2(_03653_ ), .ZN(_01287_ ) );
OAI21_X1 _17744_ ( .A(\u_lsu.pmem[4453] ), .B1(_09569_ ), .B2(_03642_ ), .ZN(_03654_ ) );
NAND3_X1 _17745_ ( .A1(_10728_ ), .A2(_09574_ ), .A3(_03550_ ), .ZN(_03655_ ) );
AOI21_X1 _17746_ ( .A(fanout_net_45 ), .B1(_03654_ ), .B2(_03655_ ), .ZN(_01288_ ) );
OAI21_X1 _17747_ ( .A(\u_lsu.pmem[4452] ), .B1(_09561_ ), .B2(_03642_ ), .ZN(_03656_ ) );
NAND3_X1 _17748_ ( .A1(_11152_ ), .A2(_09574_ ), .A3(_03550_ ), .ZN(_03657_ ) );
AOI21_X1 _17749_ ( .A(fanout_net_45 ), .B1(_03656_ ), .B2(_03657_ ), .ZN(_01289_ ) );
OAI21_X1 _17750_ ( .A(\u_lsu.pmem[4451] ), .B1(_09561_ ), .B2(_03642_ ), .ZN(_03658_ ) );
NAND3_X1 _17751_ ( .A1(_10733_ ), .A2(_09574_ ), .A3(_03550_ ), .ZN(_03659_ ) );
AOI21_X1 _17752_ ( .A(fanout_net_45 ), .B1(_03658_ ), .B2(_03659_ ), .ZN(_01290_ ) );
OAI21_X1 _17753_ ( .A(\u_lsu.pmem[4450] ), .B1(_09561_ ), .B2(_03642_ ), .ZN(_03660_ ) );
NAND3_X1 _17754_ ( .A1(_09612_ ), .A2(_09574_ ), .A3(_03550_ ), .ZN(_03661_ ) );
AOI21_X1 _17755_ ( .A(fanout_net_45 ), .B1(_03660_ ), .B2(_03661_ ), .ZN(_01291_ ) );
OAI21_X1 _17756_ ( .A(\u_lsu.pmem[4449] ), .B1(_09561_ ), .B2(_03642_ ), .ZN(_03662_ ) );
NAND3_X1 _17757_ ( .A1(_10738_ ), .A2(_09574_ ), .A3(_03550_ ), .ZN(_03663_ ) );
AOI21_X1 _17758_ ( .A(fanout_net_45 ), .B1(_03662_ ), .B2(_03663_ ), .ZN(_01292_ ) );
OAI21_X1 _17759_ ( .A(\u_lsu.pmem[4448] ), .B1(_09561_ ), .B2(_03642_ ), .ZN(_03664_ ) );
NAND3_X1 _17760_ ( .A1(_10741_ ), .A2(_09574_ ), .A3(_03550_ ), .ZN(_03665_ ) );
AOI21_X1 _17761_ ( .A(fanout_net_45 ), .B1(_03664_ ), .B2(_03665_ ), .ZN(_01293_ ) );
BUF_X4 _17762_ ( .A(_09675_ ), .Z(_03666_ ) );
OAI21_X1 _17763_ ( .A(\u_lsu.pmem[4423] ), .B1(_09639_ ), .B2(_03666_ ), .ZN(_03667_ ) );
NAND3_X1 _17764_ ( .A1(_11000_ ), .A2(_09643_ ), .A3(_03550_ ), .ZN(_03668_ ) );
AOI21_X1 _17765_ ( .A(fanout_net_45 ), .B1(_03667_ ), .B2(_03668_ ), .ZN(_01294_ ) );
OAI21_X1 _17766_ ( .A(\u_lsu.pmem[4422] ), .B1(_09639_ ), .B2(_03666_ ), .ZN(_03669_ ) );
NAND3_X1 _17767_ ( .A1(_10719_ ), .A2(_09643_ ), .A3(_09473_ ), .ZN(_03670_ ) );
AOI21_X1 _17768_ ( .A(fanout_net_45 ), .B1(_03669_ ), .B2(_03670_ ), .ZN(_01295_ ) );
OAI21_X1 _17769_ ( .A(\u_lsu.pmem[4421] ), .B1(_09639_ ), .B2(_03666_ ), .ZN(_03671_ ) );
NAND3_X1 _17770_ ( .A1(_10728_ ), .A2(_09643_ ), .A3(_09473_ ), .ZN(_03672_ ) );
AOI21_X1 _17771_ ( .A(fanout_net_45 ), .B1(_03671_ ), .B2(_03672_ ), .ZN(_01296_ ) );
BUF_X4 _17772_ ( .A(_10063_ ), .Z(_03673_ ) );
BUF_X4 _17773_ ( .A(_10578_ ), .Z(_03674_ ) );
NAND4_X1 _17774_ ( .A1(_10591_ ), .A2(_09882_ ), .A3(_03673_ ), .A4(_03674_ ), .ZN(_03675_ ) );
OAI21_X1 _17775_ ( .A(\u_lsu.pmem[3584] ), .B1(_10563_ ), .B2(_10910_ ), .ZN(_03676_ ) );
AOI21_X1 _17776_ ( .A(fanout_net_45 ), .B1(_03675_ ), .B2(_03676_ ), .ZN(_01297_ ) );
OAI21_X1 _17777_ ( .A(\u_lsu.pmem[4420] ), .B1(_09634_ ), .B2(_03666_ ), .ZN(_03677_ ) );
NAND3_X1 _17778_ ( .A1(_09589_ ), .A2(_09643_ ), .A3(_09473_ ), .ZN(_03678_ ) );
AOI21_X1 _17779_ ( .A(fanout_net_45 ), .B1(_03677_ ), .B2(_03678_ ), .ZN(_01298_ ) );
OAI21_X1 _17780_ ( .A(\u_lsu.pmem[4419] ), .B1(_09634_ ), .B2(_03666_ ), .ZN(_03679_ ) );
NAND3_X1 _17781_ ( .A1(_10733_ ), .A2(_09643_ ), .A3(_09473_ ), .ZN(_03680_ ) );
AOI21_X1 _17782_ ( .A(fanout_net_45 ), .B1(_03679_ ), .B2(_03680_ ), .ZN(_01299_ ) );
OAI21_X1 _17783_ ( .A(\u_lsu.pmem[4418] ), .B1(_09634_ ), .B2(_03666_ ), .ZN(_03681_ ) );
NAND3_X1 _17784_ ( .A1(_09612_ ), .A2(_09643_ ), .A3(_09473_ ), .ZN(_03682_ ) );
AOI21_X1 _17785_ ( .A(fanout_net_45 ), .B1(_03681_ ), .B2(_03682_ ), .ZN(_01300_ ) );
OAI21_X1 _17786_ ( .A(\u_lsu.pmem[4417] ), .B1(_09634_ ), .B2(_03666_ ), .ZN(_03683_ ) );
NAND3_X1 _17787_ ( .A1(_10738_ ), .A2(_09643_ ), .A3(_09473_ ), .ZN(_03684_ ) );
AOI21_X1 _17788_ ( .A(fanout_net_45 ), .B1(_03683_ ), .B2(_03684_ ), .ZN(_01301_ ) );
OAI21_X1 _17789_ ( .A(\u_lsu.pmem[4416] ), .B1(_09634_ ), .B2(_03666_ ), .ZN(_03685_ ) );
NAND3_X1 _17790_ ( .A1(_10741_ ), .A2(_09643_ ), .A3(_09473_ ), .ZN(_03686_ ) );
AOI21_X1 _17791_ ( .A(fanout_net_46 ), .B1(_03685_ ), .B2(_03686_ ), .ZN(_01302_ ) );
NAND4_X1 _17792_ ( .A1(_09670_ ), .A2(_03619_ ), .A3(_03622_ ), .A4(_03616_ ), .ZN(_03687_ ) );
OAI21_X1 _17793_ ( .A(\u_lsu.pmem[4391] ), .B1(_09440_ ), .B2(_09516_ ), .ZN(_03688_ ) );
AOI21_X1 _17794_ ( .A(fanout_net_46 ), .B1(_03687_ ), .B2(_03688_ ), .ZN(_01303_ ) );
NAND4_X1 _17795_ ( .A1(_09681_ ), .A2(_03619_ ), .A3(_03622_ ), .A4(_03616_ ), .ZN(_03689_ ) );
OAI21_X1 _17796_ ( .A(\u_lsu.pmem[4390] ), .B1(_09440_ ), .B2(_09516_ ), .ZN(_03690_ ) );
AOI21_X1 _17797_ ( .A(fanout_net_46 ), .B1(_03689_ ), .B2(_03690_ ), .ZN(_01304_ ) );
NAND4_X1 _17798_ ( .A1(_09685_ ), .A2(_03619_ ), .A3(_03622_ ), .A4(_03616_ ), .ZN(_03691_ ) );
OAI21_X1 _17799_ ( .A(\u_lsu.pmem[4389] ), .B1(_09440_ ), .B2(_09516_ ), .ZN(_03692_ ) );
AOI21_X1 _17800_ ( .A(fanout_net_46 ), .B1(_03691_ ), .B2(_03692_ ), .ZN(_01305_ ) );
NOR2_X1 _17801_ ( .A1(_10720_ ), .A2(_10597_ ), .ZN(_03693_ ) );
NOR2_X1 _17802_ ( .A1(_03693_ ), .A2(\u_lsu.pmem[3559] ), .ZN(_03694_ ) );
AOI211_X1 _17803_ ( .A(fanout_net_46 ), .B(_03694_ ), .C1(_09568_ ), .C2(_03693_ ), .ZN(_01306_ ) );
NAND4_X1 _17804_ ( .A1(_10603_ ), .A2(_03133_ ), .A3(_03299_ ), .A4(_03233_ ), .ZN(_03695_ ) );
OAI21_X1 _17805_ ( .A(\u_lsu.pmem[3558] ), .B1(_03205_ ), .B2(_10598_ ), .ZN(_03696_ ) );
AOI21_X1 _17806_ ( .A(fanout_net_46 ), .B1(_03695_ ), .B2(_03696_ ), .ZN(_01307_ ) );
NAND4_X1 _17807_ ( .A1(_10608_ ), .A2(_02976_ ), .A3(_03299_ ), .A4(_03233_ ), .ZN(_03697_ ) );
BUF_X4 _17808_ ( .A(_09562_ ), .Z(_03698_ ) );
OAI21_X1 _17809_ ( .A(\u_lsu.pmem[3557] ), .B1(_03698_ ), .B2(_10598_ ), .ZN(_03699_ ) );
AOI21_X1 _17810_ ( .A(fanout_net_46 ), .B1(_03697_ ), .B2(_03699_ ), .ZN(_01308_ ) );
BUF_X4 _17811_ ( .A(_10287_ ), .Z(_03700_ ) );
NAND4_X1 _17812_ ( .A1(_10611_ ), .A2(_03700_ ), .A3(_03299_ ), .A4(_03233_ ), .ZN(_03701_ ) );
OAI21_X1 _17813_ ( .A(\u_lsu.pmem[3556] ), .B1(_03698_ ), .B2(_10597_ ), .ZN(_03702_ ) );
AOI21_X1 _17814_ ( .A(fanout_net_46 ), .B1(_03701_ ), .B2(_03702_ ), .ZN(_01309_ ) );
NAND4_X1 _17815_ ( .A1(_10614_ ), .A2(_03700_ ), .A3(_03299_ ), .A4(_03233_ ), .ZN(_03703_ ) );
OAI21_X1 _17816_ ( .A(\u_lsu.pmem[3555] ), .B1(_03698_ ), .B2(_10597_ ), .ZN(_03704_ ) );
AOI21_X1 _17817_ ( .A(fanout_net_46 ), .B1(_03703_ ), .B2(_03704_ ), .ZN(_01310_ ) );
BUF_X4 _17818_ ( .A(_09459_ ), .Z(_03705_ ) );
OAI21_X1 _17819_ ( .A(\u_lsu.pmem[4295] ), .B1(_03705_ ), .B2(_09808_ ), .ZN(_03706_ ) );
NAND4_X1 _17820_ ( .A1(_09742_ ), .A2(_03504_ ), .A3(_03640_ ), .A4(_09798_ ), .ZN(_03707_ ) );
AOI21_X1 _17821_ ( .A(fanout_net_46 ), .B1(_03706_ ), .B2(_03707_ ), .ZN(_01311_ ) );
NAND4_X1 _17822_ ( .A1(_10617_ ), .A2(_03700_ ), .A3(_03299_ ), .A4(_03233_ ), .ZN(_03708_ ) );
OAI21_X1 _17823_ ( .A(\u_lsu.pmem[3554] ), .B1(_03698_ ), .B2(_10597_ ), .ZN(_03709_ ) );
AOI21_X1 _17824_ ( .A(fanout_net_46 ), .B1(_03708_ ), .B2(_03709_ ), .ZN(_01312_ ) );
BUF_X4 _17825_ ( .A(_11492_ ), .Z(_03710_ ) );
NAND4_X1 _17826_ ( .A1(_10621_ ), .A2(_03133_ ), .A3(_03299_ ), .A4(_03710_ ), .ZN(_03711_ ) );
OAI21_X1 _17827_ ( .A(\u_lsu.pmem[3553] ), .B1(_03698_ ), .B2(_10597_ ), .ZN(_03712_ ) );
AOI21_X1 _17828_ ( .A(fanout_net_46 ), .B1(_03711_ ), .B2(_03712_ ), .ZN(_01313_ ) );
NAND4_X1 _17829_ ( .A1(_10624_ ), .A2(_03700_ ), .A3(_03299_ ), .A4(_03710_ ), .ZN(_03713_ ) );
OAI21_X1 _17830_ ( .A(\u_lsu.pmem[3552] ), .B1(_03698_ ), .B2(_10597_ ), .ZN(_03714_ ) );
AOI21_X1 _17831_ ( .A(fanout_net_46 ), .B1(_03713_ ), .B2(_03714_ ), .ZN(_01314_ ) );
NOR2_X1 _17832_ ( .A1(_10720_ ), .A2(_10628_ ), .ZN(_03715_ ) );
NOR2_X1 _17833_ ( .A1(_03715_ ), .A2(\u_lsu.pmem[3527] ), .ZN(_03716_ ) );
AOI211_X1 _17834_ ( .A(fanout_net_46 ), .B(_03716_ ), .C1(_09568_ ), .C2(_03715_ ), .ZN(_01315_ ) );
BUF_X4 _17835_ ( .A(_02196_ ), .Z(_03717_ ) );
NAND4_X1 _17836_ ( .A1(_10632_ ), .A2(_03700_ ), .A3(_03717_ ), .A4(_03710_ ), .ZN(_03718_ ) );
OAI21_X1 _17837_ ( .A(\u_lsu.pmem[3526] ), .B1(_03698_ ), .B2(_10629_ ), .ZN(_03719_ ) );
AOI21_X1 _17838_ ( .A(fanout_net_46 ), .B1(_03718_ ), .B2(_03719_ ), .ZN(_01316_ ) );
NAND4_X1 _17839_ ( .A1(_10635_ ), .A2(_03700_ ), .A3(_03717_ ), .A4(_03710_ ), .ZN(_03720_ ) );
OAI21_X1 _17840_ ( .A(\u_lsu.pmem[3525] ), .B1(_03698_ ), .B2(_10629_ ), .ZN(_03721_ ) );
AOI21_X1 _17841_ ( .A(fanout_net_46 ), .B1(_03720_ ), .B2(_03721_ ), .ZN(_01317_ ) );
NAND4_X1 _17842_ ( .A1(_10641_ ), .A2(_03700_ ), .A3(_03717_ ), .A4(_03710_ ), .ZN(_03722_ ) );
OAI21_X1 _17843_ ( .A(\u_lsu.pmem[3524] ), .B1(_03698_ ), .B2(_10628_ ), .ZN(_03723_ ) );
AOI21_X1 _17844_ ( .A(fanout_net_46 ), .B1(_03722_ ), .B2(_03723_ ), .ZN(_01318_ ) );
NAND4_X1 _17845_ ( .A1(_10645_ ), .A2(_03700_ ), .A3(_03717_ ), .A4(_03710_ ), .ZN(_03724_ ) );
OAI21_X1 _17846_ ( .A(\u_lsu.pmem[3523] ), .B1(_03698_ ), .B2(_10628_ ), .ZN(_03725_ ) );
AOI21_X1 _17847_ ( .A(fanout_net_46 ), .B1(_03724_ ), .B2(_03725_ ), .ZN(_01319_ ) );
NAND4_X1 _17848_ ( .A1(_10649_ ), .A2(_03700_ ), .A3(_03717_ ), .A4(_03710_ ), .ZN(_03726_ ) );
BUF_X4 _17849_ ( .A(_09562_ ), .Z(_03727_ ) );
OAI21_X1 _17850_ ( .A(\u_lsu.pmem[3522] ), .B1(_03727_ ), .B2(_10628_ ), .ZN(_03728_ ) );
AOI21_X1 _17851_ ( .A(fanout_net_46 ), .B1(_03726_ ), .B2(_03728_ ), .ZN(_01320_ ) );
NAND4_X1 _17852_ ( .A1(_10652_ ), .A2(_03133_ ), .A3(_03717_ ), .A4(_03710_ ), .ZN(_03729_ ) );
OAI21_X1 _17853_ ( .A(\u_lsu.pmem[3521] ), .B1(_03727_ ), .B2(_10628_ ), .ZN(_03730_ ) );
AOI21_X1 _17854_ ( .A(fanout_net_46 ), .B1(_03729_ ), .B2(_03730_ ), .ZN(_01321_ ) );
NAND4_X1 _17855_ ( .A1(_09804_ ), .A2(_09806_ ), .A3(_03622_ ), .A4(_03616_ ), .ZN(_03731_ ) );
OAI21_X1 _17856_ ( .A(\u_lsu.pmem[4294] ), .B1(_03606_ ), .B2(_09808_ ), .ZN(_03732_ ) );
AOI21_X1 _17857_ ( .A(fanout_net_46 ), .B1(_03731_ ), .B2(_03732_ ), .ZN(_01322_ ) );
NAND4_X1 _17858_ ( .A1(_10655_ ), .A2(_03700_ ), .A3(_03717_ ), .A4(_03710_ ), .ZN(_03733_ ) );
OAI21_X1 _17859_ ( .A(\u_lsu.pmem[3520] ), .B1(_03727_ ), .B2(_10628_ ), .ZN(_03734_ ) );
AOI21_X1 _17860_ ( .A(fanout_net_46 ), .B1(_03733_ ), .B2(_03734_ ), .ZN(_01323_ ) );
BUF_X4 _17861_ ( .A(_10287_ ), .Z(_03735_ ) );
NAND4_X1 _17862_ ( .A1(_10658_ ), .A2(_03735_ ), .A3(_03717_ ), .A4(_03710_ ), .ZN(_03736_ ) );
OAI21_X1 _17863_ ( .A(\u_lsu.pmem[3495] ), .B1(_03727_ ), .B2(_10663_ ), .ZN(_03737_ ) );
AOI21_X1 _17864_ ( .A(fanout_net_46 ), .B1(_03736_ ), .B2(_03737_ ), .ZN(_01324_ ) );
BUF_X4 _17865_ ( .A(_11492_ ), .Z(_03738_ ) );
NAND4_X1 _17866_ ( .A1(_10665_ ), .A2(_03133_ ), .A3(_03717_ ), .A4(_03738_ ), .ZN(_03739_ ) );
OAI21_X1 _17867_ ( .A(\u_lsu.pmem[3494] ), .B1(_03727_ ), .B2(_10663_ ), .ZN(_03740_ ) );
AOI21_X1 _17868_ ( .A(fanout_net_46 ), .B1(_03739_ ), .B2(_03740_ ), .ZN(_01325_ ) );
NAND4_X1 _17869_ ( .A1(_10668_ ), .A2(_03735_ ), .A3(_03717_ ), .A4(_03738_ ), .ZN(_03741_ ) );
OAI21_X1 _17870_ ( .A(\u_lsu.pmem[3493] ), .B1(_03727_ ), .B2(_10662_ ), .ZN(_03742_ ) );
AOI21_X1 _17871_ ( .A(fanout_net_46 ), .B1(_03741_ ), .B2(_03742_ ), .ZN(_01326_ ) );
BUF_X4 _17872_ ( .A(_03020_ ), .Z(_03743_ ) );
BUF_X4 _17873_ ( .A(_02196_ ), .Z(_03744_ ) );
NAND4_X1 _17874_ ( .A1(_10671_ ), .A2(_03743_ ), .A3(_03744_ ), .A4(_03738_ ), .ZN(_03745_ ) );
OAI21_X1 _17875_ ( .A(\u_lsu.pmem[3492] ), .B1(_03727_ ), .B2(_10662_ ), .ZN(_03746_ ) );
AOI21_X1 _17876_ ( .A(fanout_net_46 ), .B1(_03745_ ), .B2(_03746_ ), .ZN(_01327_ ) );
NAND4_X1 _17877_ ( .A1(_10674_ ), .A2(_03743_ ), .A3(_03744_ ), .A4(_03738_ ), .ZN(_03747_ ) );
OAI21_X1 _17878_ ( .A(\u_lsu.pmem[3491] ), .B1(_03727_ ), .B2(_10662_ ), .ZN(_03748_ ) );
AOI21_X1 _17879_ ( .A(fanout_net_46 ), .B1(_03747_ ), .B2(_03748_ ), .ZN(_01328_ ) );
NAND4_X1 _17880_ ( .A1(_10679_ ), .A2(_03743_ ), .A3(_03744_ ), .A4(_03738_ ), .ZN(_03749_ ) );
OAI21_X1 _17881_ ( .A(\u_lsu.pmem[3490] ), .B1(_03727_ ), .B2(_10662_ ), .ZN(_03750_ ) );
AOI21_X1 _17882_ ( .A(fanout_net_46 ), .B1(_03749_ ), .B2(_03750_ ), .ZN(_01329_ ) );
NAND4_X1 _17883_ ( .A1(_10682_ ), .A2(_03743_ ), .A3(_03744_ ), .A4(_03738_ ), .ZN(_03751_ ) );
OAI21_X1 _17884_ ( .A(\u_lsu.pmem[3489] ), .B1(_03727_ ), .B2(_10662_ ), .ZN(_03752_ ) );
AOI21_X1 _17885_ ( .A(fanout_net_46 ), .B1(_03751_ ), .B2(_03752_ ), .ZN(_01330_ ) );
BUF_X4 _17886_ ( .A(_09621_ ), .Z(_03753_ ) );
NAND4_X1 _17887_ ( .A1(_02903_ ), .A2(_02935_ ), .A3(_03753_ ), .A4(_10661_ ), .ZN(_03754_ ) );
BUF_X4 _17888_ ( .A(_09562_ ), .Z(_03755_ ) );
OAI21_X1 _17889_ ( .A(\u_lsu.pmem[3488] ), .B1(_03755_ ), .B2(_10662_ ), .ZN(_03756_ ) );
AOI21_X1 _17890_ ( .A(fanout_net_46 ), .B1(_03754_ ), .B2(_03756_ ), .ZN(_01331_ ) );
OAI21_X1 _17891_ ( .A(\u_lsu.pmem[3463] ), .B1(_10692_ ), .B2(_09911_ ), .ZN(_03757_ ) );
NAND4_X1 _17892_ ( .A1(_02869_ ), .A2(_03478_ ), .A3(_02672_ ), .A4(_02526_ ), .ZN(_03758_ ) );
AOI21_X1 _17893_ ( .A(fanout_net_47 ), .B1(_03757_ ), .B2(_03758_ ), .ZN(_01332_ ) );
NAND4_X1 _17894_ ( .A1(_09811_ ), .A2(_03619_ ), .A3(_03622_ ), .A4(_03616_ ), .ZN(_03759_ ) );
OAI21_X1 _17895_ ( .A(\u_lsu.pmem[4293] ), .B1(_03606_ ), .B2(_09808_ ), .ZN(_03760_ ) );
AOI21_X1 _17896_ ( .A(fanout_net_47 ), .B1(_03759_ ), .B2(_03760_ ), .ZN(_01333_ ) );
OAI21_X1 _17897_ ( .A(\u_lsu.pmem[3462] ), .B1(_10692_ ), .B2(_09911_ ), .ZN(_03761_ ) );
NAND4_X1 _17898_ ( .A1(_02869_ ), .A2(_03056_ ), .A3(_02672_ ), .A4(_02526_ ), .ZN(_03762_ ) );
AOI21_X1 _17899_ ( .A(fanout_net_47 ), .B1(_03761_ ), .B2(_03762_ ), .ZN(_01334_ ) );
OAI21_X1 _17900_ ( .A(\u_lsu.pmem[3461] ), .B1(_10691_ ), .B2(_09911_ ), .ZN(_03763_ ) );
NAND4_X1 _17901_ ( .A1(_02869_ ), .A2(_03059_ ), .A3(_02672_ ), .A4(_02526_ ), .ZN(_03764_ ) );
AOI21_X1 _17902_ ( .A(fanout_net_47 ), .B1(_03763_ ), .B2(_03764_ ), .ZN(_01335_ ) );
OAI21_X1 _17903_ ( .A(\u_lsu.pmem[3460] ), .B1(_10691_ ), .B2(_09911_ ), .ZN(_03765_ ) );
NAND4_X1 _17904_ ( .A1(_02869_ ), .A2(_03064_ ), .A3(_02672_ ), .A4(_02526_ ), .ZN(_03766_ ) );
AOI21_X1 _17905_ ( .A(fanout_net_47 ), .B1(_03765_ ), .B2(_03766_ ), .ZN(_01336_ ) );
OAI21_X1 _17906_ ( .A(\u_lsu.pmem[3459] ), .B1(_10691_ ), .B2(_09911_ ), .ZN(_03767_ ) );
NAND4_X1 _17907_ ( .A1(_02869_ ), .A2(_10915_ ), .A3(_02672_ ), .A4(_02526_ ), .ZN(_03768_ ) );
AOI21_X1 _17908_ ( .A(fanout_net_47 ), .B1(_03767_ ), .B2(_03768_ ), .ZN(_01337_ ) );
BUF_X4 _17909_ ( .A(_09647_ ), .Z(_03769_ ) );
OAI21_X1 _17910_ ( .A(\u_lsu.pmem[3458] ), .B1(_10691_ ), .B2(_03769_ ), .ZN(_03770_ ) );
NAND4_X1 _17911_ ( .A1(_09537_ ), .A2(_03107_ ), .A3(_02672_ ), .A4(_02526_ ), .ZN(_03771_ ) );
AOI21_X1 _17912_ ( .A(fanout_net_47 ), .B1(_03770_ ), .B2(_03771_ ), .ZN(_01338_ ) );
OAI21_X1 _17913_ ( .A(\u_lsu.pmem[3457] ), .B1(_10691_ ), .B2(_03769_ ), .ZN(_03772_ ) );
NAND4_X1 _17914_ ( .A1(_02869_ ), .A2(_02308_ ), .A3(_02672_ ), .A4(_02526_ ), .ZN(_03773_ ) );
AOI21_X1 _17915_ ( .A(fanout_net_47 ), .B1(_03772_ ), .B2(_03773_ ), .ZN(_01339_ ) );
OAI21_X1 _17916_ ( .A(\u_lsu.pmem[3456] ), .B1(_10691_ ), .B2(_03769_ ), .ZN(_03774_ ) );
NAND4_X1 _17917_ ( .A1(_10694_ ), .A2(_11131_ ), .A3(_02672_ ), .A4(_02526_ ), .ZN(_03775_ ) );
AOI21_X1 _17918_ ( .A(fanout_net_47 ), .B1(_03774_ ), .B2(_03775_ ), .ZN(_01340_ ) );
NOR2_X1 _17919_ ( .A1(_10716_ ), .A2(_10046_ ), .ZN(_03776_ ) );
OAI21_X1 _17920_ ( .A(_10715_ ), .B1(_03776_ ), .B2(\u_lsu.pmem[3431] ), .ZN(_03777_ ) );
AOI21_X1 _17921_ ( .A(_03777_ ), .B1(_09638_ ), .B2(_03776_ ), .ZN(_01341_ ) );
NAND4_X1 _17922_ ( .A1(_02903_ ), .A2(_09925_ ), .A3(_03744_ ), .A4(_10724_ ), .ZN(_03778_ ) );
OAI21_X1 _17923_ ( .A(\u_lsu.pmem[3430] ), .B1(_10726_ ), .B2(_10910_ ), .ZN(_03779_ ) );
AOI21_X1 _17924_ ( .A(fanout_net_47 ), .B1(_03778_ ), .B2(_03779_ ), .ZN(_01342_ ) );
NAND4_X1 _17925_ ( .A1(_02903_ ), .A2(_09928_ ), .A3(_03744_ ), .A4(_10724_ ), .ZN(_03780_ ) );
OAI21_X1 _17926_ ( .A(\u_lsu.pmem[3429] ), .B1(_10726_ ), .B2(_10910_ ), .ZN(_03781_ ) );
AOI21_X1 _17927_ ( .A(fanout_net_47 ), .B1(_03780_ ), .B2(_03781_ ), .ZN(_01343_ ) );
NAND4_X1 _17928_ ( .A1(_09815_ ), .A2(_03619_ ), .A3(_03622_ ), .A4(_03616_ ), .ZN(_03782_ ) );
OAI21_X1 _17929_ ( .A(\u_lsu.pmem[4292] ), .B1(_03606_ ), .B2(_09799_ ), .ZN(_03783_ ) );
AOI21_X1 _17930_ ( .A(fanout_net_47 ), .B1(_03782_ ), .B2(_03783_ ), .ZN(_01344_ ) );
NAND4_X1 _17931_ ( .A1(_02903_ ), .A2(_09931_ ), .A3(_03744_ ), .A4(_10724_ ), .ZN(_03784_ ) );
OAI21_X1 _17932_ ( .A(\u_lsu.pmem[3428] ), .B1(_10726_ ), .B2(_10910_ ), .ZN(_03785_ ) );
AOI21_X1 _17933_ ( .A(fanout_net_47 ), .B1(_03784_ ), .B2(_03785_ ), .ZN(_01345_ ) );
BUF_X4 _17934_ ( .A(_10723_ ), .Z(_03786_ ) );
NAND4_X1 _17935_ ( .A1(_02903_ ), .A2(_03091_ ), .A3(_03744_ ), .A4(_03786_ ), .ZN(_03787_ ) );
OAI21_X1 _17936_ ( .A(\u_lsu.pmem[3427] ), .B1(_10726_ ), .B2(_10910_ ), .ZN(_03788_ ) );
AOI21_X1 _17937_ ( .A(fanout_net_47 ), .B1(_03787_ ), .B2(_03788_ ), .ZN(_01346_ ) );
NAND4_X1 _17938_ ( .A1(_02903_ ), .A2(_09938_ ), .A3(_03744_ ), .A4(_03786_ ), .ZN(_03789_ ) );
OAI21_X1 _17939_ ( .A(\u_lsu.pmem[3426] ), .B1(_10726_ ), .B2(_10910_ ), .ZN(_03790_ ) );
AOI21_X1 _17940_ ( .A(fanout_net_47 ), .B1(_03789_ ), .B2(_03790_ ), .ZN(_01347_ ) );
NAND4_X1 _17941_ ( .A1(_02903_ ), .A2(_03143_ ), .A3(_03744_ ), .A4(_03786_ ), .ZN(_03791_ ) );
OAI21_X1 _17942_ ( .A(\u_lsu.pmem[3425] ), .B1(_10726_ ), .B2(_10910_ ), .ZN(_03792_ ) );
AOI21_X1 _17943_ ( .A(fanout_net_47 ), .B1(_03791_ ), .B2(_03792_ ), .ZN(_01348_ ) );
BUF_X4 _17944_ ( .A(_09953_ ), .Z(_03793_ ) );
BUF_X4 _17945_ ( .A(_02196_ ), .Z(_03794_ ) );
NAND4_X1 _17946_ ( .A1(_03793_ ), .A2(_09944_ ), .A3(_03794_ ), .A4(_03786_ ), .ZN(_03795_ ) );
BUF_X4 _17947_ ( .A(_10046_ ), .Z(_03796_ ) );
OAI21_X1 _17948_ ( .A(\u_lsu.pmem[3424] ), .B1(_10726_ ), .B2(_03796_ ), .ZN(_03797_ ) );
AOI21_X1 _17949_ ( .A(fanout_net_47 ), .B1(_03795_ ), .B2(_03797_ ), .ZN(_01349_ ) );
AND2_X1 _17950_ ( .A1(_10746_ ), .A2(_10012_ ), .ZN(_03798_ ) );
OAI21_X1 _17951_ ( .A(_10715_ ), .B1(_03798_ ), .B2(\u_lsu.pmem[3399] ), .ZN(_03799_ ) );
AOI21_X1 _17952_ ( .A(_03799_ ), .B1(_09638_ ), .B2(_03798_ ), .ZN(_01350_ ) );
NAND4_X1 _17953_ ( .A1(_03793_ ), .A2(_09925_ ), .A3(_03794_ ), .A4(_10751_ ), .ZN(_03800_ ) );
OAI21_X1 _17954_ ( .A(\u_lsu.pmem[3398] ), .B1(_10748_ ), .B2(_03796_ ), .ZN(_03801_ ) );
AOI21_X1 _17955_ ( .A(fanout_net_47 ), .B1(_03800_ ), .B2(_03801_ ), .ZN(_01351_ ) );
NAND4_X1 _17956_ ( .A1(_03793_ ), .A2(_09928_ ), .A3(_03794_ ), .A4(_10751_ ), .ZN(_03802_ ) );
OAI21_X1 _17957_ ( .A(\u_lsu.pmem[3397] ), .B1(_10748_ ), .B2(_03796_ ), .ZN(_03803_ ) );
AOI21_X1 _17958_ ( .A(fanout_net_47 ), .B1(_03802_ ), .B2(_03803_ ), .ZN(_01352_ ) );
BUF_X4 _17959_ ( .A(_10745_ ), .Z(_03804_ ) );
NAND4_X1 _17960_ ( .A1(_03793_ ), .A2(_09931_ ), .A3(_03794_ ), .A4(_03804_ ), .ZN(_03805_ ) );
OAI21_X1 _17961_ ( .A(\u_lsu.pmem[3396] ), .B1(_10747_ ), .B2(_03796_ ), .ZN(_03806_ ) );
AOI21_X1 _17962_ ( .A(fanout_net_47 ), .B1(_03805_ ), .B2(_03806_ ), .ZN(_01353_ ) );
NAND4_X1 _17963_ ( .A1(_03793_ ), .A2(_03091_ ), .A3(_03794_ ), .A4(_03804_ ), .ZN(_03807_ ) );
OAI21_X1 _17964_ ( .A(\u_lsu.pmem[3395] ), .B1(_10747_ ), .B2(_03796_ ), .ZN(_03808_ ) );
AOI21_X1 _17965_ ( .A(fanout_net_47 ), .B1(_03807_ ), .B2(_03808_ ), .ZN(_01354_ ) );
NAND4_X1 _17966_ ( .A1(_09819_ ), .A2(_03619_ ), .A3(_03622_ ), .A4(_03616_ ), .ZN(_03809_ ) );
BUF_X4 _17967_ ( .A(_09443_ ), .Z(_03810_ ) );
OAI21_X1 _17968_ ( .A(\u_lsu.pmem[4291] ), .B1(_03810_ ), .B2(_09799_ ), .ZN(_03811_ ) );
AOI21_X1 _17969_ ( .A(fanout_net_47 ), .B1(_03809_ ), .B2(_03811_ ), .ZN(_01355_ ) );
NAND4_X1 _17970_ ( .A1(_03793_ ), .A2(_09938_ ), .A3(_03794_ ), .A4(_03804_ ), .ZN(_03812_ ) );
OAI21_X1 _17971_ ( .A(\u_lsu.pmem[3394] ), .B1(_10747_ ), .B2(_03796_ ), .ZN(_03813_ ) );
AOI21_X1 _17972_ ( .A(fanout_net_47 ), .B1(_03812_ ), .B2(_03813_ ), .ZN(_01356_ ) );
NAND4_X1 _17973_ ( .A1(_03793_ ), .A2(_03143_ ), .A3(_03794_ ), .A4(_03804_ ), .ZN(_03814_ ) );
OAI21_X1 _17974_ ( .A(\u_lsu.pmem[3393] ), .B1(_10747_ ), .B2(_03796_ ), .ZN(_03815_ ) );
AOI21_X1 _17975_ ( .A(fanout_net_47 ), .B1(_03814_ ), .B2(_03815_ ), .ZN(_01357_ ) );
NAND4_X1 _17976_ ( .A1(_03793_ ), .A2(_09944_ ), .A3(_03794_ ), .A4(_03804_ ), .ZN(_03816_ ) );
OAI21_X1 _17977_ ( .A(\u_lsu.pmem[3392] ), .B1(_10747_ ), .B2(_03796_ ), .ZN(_03817_ ) );
AOI21_X1 _17978_ ( .A(fanout_net_47 ), .B1(_03816_ ), .B2(_03817_ ), .ZN(_01358_ ) );
NAND4_X1 _17979_ ( .A1(_09670_ ), .A2(_03743_ ), .A3(_03794_ ), .A4(_03738_ ), .ZN(_03818_ ) );
OAI21_X1 _17980_ ( .A(\u_lsu.pmem[3367] ), .B1(_10775_ ), .B2(_02584_ ), .ZN(_03819_ ) );
AOI21_X1 _17981_ ( .A(fanout_net_47 ), .B1(_03818_ ), .B2(_03819_ ), .ZN(_01359_ ) );
NAND4_X1 _17982_ ( .A1(_09681_ ), .A2(_03743_ ), .A3(_03794_ ), .A4(_03738_ ), .ZN(_03820_ ) );
OAI21_X1 _17983_ ( .A(\u_lsu.pmem[3366] ), .B1(_10775_ ), .B2(_02584_ ), .ZN(_03821_ ) );
AOI21_X1 _17984_ ( .A(fanout_net_47 ), .B1(_03820_ ), .B2(_03821_ ), .ZN(_01360_ ) );
BUF_X4 _17985_ ( .A(_02196_ ), .Z(_03822_ ) );
NAND4_X1 _17986_ ( .A1(_09685_ ), .A2(_03743_ ), .A3(_03822_ ), .A4(_03738_ ), .ZN(_03823_ ) );
OAI21_X1 _17987_ ( .A(\u_lsu.pmem[3365] ), .B1(_10775_ ), .B2(_02584_ ), .ZN(_03824_ ) );
AOI21_X1 _17988_ ( .A(fanout_net_47 ), .B1(_03823_ ), .B2(_03824_ ), .ZN(_01361_ ) );
OAI21_X1 _17989_ ( .A(\u_lsu.pmem[3364] ), .B1(_10776_ ), .B2(_03769_ ), .ZN(_03825_ ) );
BUF_X4 _17990_ ( .A(_09641_ ), .Z(_03826_ ) );
NAND3_X1 _17991_ ( .A1(_03826_ ), .A2(_09589_ ), .A3(_10774_ ), .ZN(_03827_ ) );
AOI21_X1 _17992_ ( .A(fanout_net_47 ), .B1(_03825_ ), .B2(_03827_ ), .ZN(_01362_ ) );
OAI21_X1 _17993_ ( .A(\u_lsu.pmem[3363] ), .B1(_10776_ ), .B2(_03769_ ), .ZN(_03828_ ) );
NAND3_X1 _17994_ ( .A1(_03826_ ), .A2(_09592_ ), .A3(_10774_ ), .ZN(_03829_ ) );
AOI21_X1 _17995_ ( .A(fanout_net_47 ), .B1(_03828_ ), .B2(_03829_ ), .ZN(_01363_ ) );
OAI21_X1 _17996_ ( .A(\u_lsu.pmem[3362] ), .B1(_10776_ ), .B2(_03769_ ), .ZN(_03830_ ) );
NAND3_X1 _17997_ ( .A1(_03826_ ), .A2(_09695_ ), .A3(_10774_ ), .ZN(_03831_ ) );
AOI21_X1 _17998_ ( .A(fanout_net_48 ), .B1(_03830_ ), .B2(_03831_ ), .ZN(_01364_ ) );
OAI21_X1 _17999_ ( .A(\u_lsu.pmem[3361] ), .B1(_10776_ ), .B2(_03769_ ), .ZN(_03832_ ) );
NAND3_X1 _18000_ ( .A1(_03826_ ), .A2(_09617_ ), .A3(_10774_ ), .ZN(_03833_ ) );
AOI21_X1 _18001_ ( .A(fanout_net_48 ), .B1(_03832_ ), .B2(_03833_ ), .ZN(_01365_ ) );
BUF_X4 _18002_ ( .A(_09730_ ), .Z(_03834_ ) );
NAND4_X1 _18003_ ( .A1(_09827_ ), .A2(_03619_ ), .A3(_03622_ ), .A4(_03834_ ), .ZN(_03835_ ) );
OAI21_X1 _18004_ ( .A(\u_lsu.pmem[4290] ), .B1(_03810_ ), .B2(_09799_ ), .ZN(_03836_ ) );
AOI21_X1 _18005_ ( .A(fanout_net_48 ), .B1(_03835_ ), .B2(_03836_ ), .ZN(_01366_ ) );
NAND4_X1 _18006_ ( .A1(_09703_ ), .A2(_03743_ ), .A3(_03822_ ), .A4(_03738_ ), .ZN(_03837_ ) );
OAI21_X1 _18007_ ( .A(\u_lsu.pmem[3360] ), .B1(_10775_ ), .B2(_02584_ ), .ZN(_03838_ ) );
AOI21_X1 _18008_ ( .A(fanout_net_48 ), .B1(_03837_ ), .B2(_03838_ ), .ZN(_01367_ ) );
BUF_X4 _18009_ ( .A(_11492_ ), .Z(_03839_ ) );
NAND4_X1 _18010_ ( .A1(_09708_ ), .A2(_03735_ ), .A3(_03822_ ), .A4(_03839_ ), .ZN(_03840_ ) );
OAI21_X1 _18011_ ( .A(\u_lsu.pmem[3335] ), .B1(_03755_ ), .B2(_10799_ ), .ZN(_03841_ ) );
AOI21_X1 _18012_ ( .A(fanout_net_48 ), .B1(_03840_ ), .B2(_03841_ ), .ZN(_01368_ ) );
NAND4_X1 _18013_ ( .A1(_09715_ ), .A2(_10974_ ), .A3(_10876_ ), .A4(_03674_ ), .ZN(_03842_ ) );
OAI21_X1 _18014_ ( .A(\u_lsu.pmem[3334] ), .B1(_03755_ ), .B2(_10799_ ), .ZN(_03843_ ) );
AOI21_X1 _18015_ ( .A(fanout_net_48 ), .B1(_03842_ ), .B2(_03843_ ), .ZN(_01369_ ) );
NAND4_X1 _18016_ ( .A1(_09718_ ), .A2(_10974_ ), .A3(_10876_ ), .A4(_03674_ ), .ZN(_03844_ ) );
OAI21_X1 _18017_ ( .A(\u_lsu.pmem[3333] ), .B1(_03755_ ), .B2(_10798_ ), .ZN(_03845_ ) );
AOI21_X1 _18018_ ( .A(fanout_net_48 ), .B1(_03844_ ), .B2(_03845_ ), .ZN(_01370_ ) );
NAND4_X1 _18019_ ( .A1(_09721_ ), .A2(_10974_ ), .A3(_10876_ ), .A4(_03674_ ), .ZN(_03846_ ) );
OAI21_X1 _18020_ ( .A(\u_lsu.pmem[3332] ), .B1(_03755_ ), .B2(_10798_ ), .ZN(_03847_ ) );
AOI21_X1 _18021_ ( .A(fanout_net_48 ), .B1(_03846_ ), .B2(_03847_ ), .ZN(_01371_ ) );
NAND4_X1 _18022_ ( .A1(_09725_ ), .A2(_10974_ ), .A3(_10876_ ), .A4(_03674_ ), .ZN(_03848_ ) );
OAI21_X1 _18023_ ( .A(\u_lsu.pmem[3331] ), .B1(_03755_ ), .B2(_10798_ ), .ZN(_03849_ ) );
AOI21_X1 _18024_ ( .A(fanout_net_48 ), .B1(_03848_ ), .B2(_03849_ ), .ZN(_01372_ ) );
BUF_X4 _18025_ ( .A(_09471_ ), .Z(_03850_ ) );
NOR2_X1 _18026_ ( .A1(_03850_ ), .A2(_10798_ ), .ZN(_03851_ ) );
NOR2_X1 _18027_ ( .A1(_03851_ ), .A2(\u_lsu.pmem[3330] ), .ZN(_03852_ ) );
AOI211_X1 _18028_ ( .A(fanout_net_48 ), .B(_03852_ ), .C1(_09973_ ), .C2(_03851_ ), .ZN(_01373_ ) );
NAND4_X1 _18029_ ( .A1(_09733_ ), .A2(_03743_ ), .A3(_03822_ ), .A4(_03839_ ), .ZN(_03853_ ) );
OAI21_X1 _18030_ ( .A(\u_lsu.pmem[3329] ), .B1(_03755_ ), .B2(_10798_ ), .ZN(_03854_ ) );
AOI21_X1 _18031_ ( .A(fanout_net_48 ), .B1(_03853_ ), .B2(_03854_ ), .ZN(_01374_ ) );
NAND4_X1 _18032_ ( .A1(_09736_ ), .A2(_10974_ ), .A3(_10876_ ), .A4(_03674_ ), .ZN(_03855_ ) );
OAI21_X1 _18033_ ( .A(\u_lsu.pmem[3328] ), .B1(_03755_ ), .B2(_10798_ ), .ZN(_03856_ ) );
AOI21_X1 _18034_ ( .A(fanout_net_48 ), .B1(_03855_ ), .B2(_03856_ ), .ZN(_01375_ ) );
NAND4_X1 _18035_ ( .A1(_03793_ ), .A2(_02935_ ), .A3(_09914_ ), .A4(_10819_ ), .ZN(_03857_ ) );
OAI21_X1 _18036_ ( .A(\u_lsu.pmem[3303] ), .B1(_03755_ ), .B2(_10821_ ), .ZN(_03858_ ) );
AOI21_X1 _18037_ ( .A(fanout_net_48 ), .B1(_03857_ ), .B2(_03858_ ), .ZN(_01376_ ) );
NAND4_X1 _18038_ ( .A1(_09831_ ), .A2(_03619_ ), .A3(_03622_ ), .A4(_03834_ ), .ZN(_03859_ ) );
OAI21_X1 _18039_ ( .A(\u_lsu.pmem[4289] ), .B1(_03810_ ), .B2(_09799_ ), .ZN(_03860_ ) );
AOI21_X1 _18040_ ( .A(fanout_net_48 ), .B1(_03859_ ), .B2(_03860_ ), .ZN(_01377_ ) );
NAND4_X1 _18041_ ( .A1(_09756_ ), .A2(_03735_ ), .A3(_03822_ ), .A4(_03839_ ), .ZN(_03861_ ) );
OAI21_X1 _18042_ ( .A(\u_lsu.pmem[3302] ), .B1(_03755_ ), .B2(_10821_ ), .ZN(_03862_ ) );
AOI21_X1 _18043_ ( .A(fanout_net_48 ), .B1(_03861_ ), .B2(_03862_ ), .ZN(_01378_ ) );
NAND4_X1 _18044_ ( .A1(_09763_ ), .A2(_03743_ ), .A3(_03822_ ), .A4(_03839_ ), .ZN(_03863_ ) );
BUF_X4 _18045_ ( .A(_09562_ ), .Z(_03864_ ) );
OAI21_X1 _18046_ ( .A(\u_lsu.pmem[3301] ), .B1(_03864_ ), .B2(_10820_ ), .ZN(_03865_ ) );
AOI21_X1 _18047_ ( .A(fanout_net_48 ), .B1(_03863_ ), .B2(_03865_ ), .ZN(_01379_ ) );
NAND4_X1 _18048_ ( .A1(_09770_ ), .A2(_03735_ ), .A3(_03822_ ), .A4(_03839_ ), .ZN(_03866_ ) );
OAI21_X1 _18049_ ( .A(\u_lsu.pmem[3300] ), .B1(_03864_ ), .B2(_10820_ ), .ZN(_03867_ ) );
AOI21_X1 _18050_ ( .A(fanout_net_48 ), .B1(_03866_ ), .B2(_03867_ ), .ZN(_01380_ ) );
BUF_X4 _18051_ ( .A(_03020_ ), .Z(_03868_ ) );
NAND4_X1 _18052_ ( .A1(_09775_ ), .A2(_03868_ ), .A3(_03822_ ), .A4(_03839_ ), .ZN(_03869_ ) );
OAI21_X1 _18053_ ( .A(\u_lsu.pmem[3299] ), .B1(_03864_ ), .B2(_10820_ ), .ZN(_03870_ ) );
AOI21_X1 _18054_ ( .A(fanout_net_48 ), .B1(_03869_ ), .B2(_03870_ ), .ZN(_01381_ ) );
NAND4_X1 _18055_ ( .A1(_09780_ ), .A2(_03868_ ), .A3(_03822_ ), .A4(_03839_ ), .ZN(_03871_ ) );
OAI21_X1 _18056_ ( .A(\u_lsu.pmem[3298] ), .B1(_03864_ ), .B2(_10820_ ), .ZN(_03872_ ) );
AOI21_X1 _18057_ ( .A(fanout_net_48 ), .B1(_03871_ ), .B2(_03872_ ), .ZN(_01382_ ) );
NAND4_X1 _18058_ ( .A1(_09787_ ), .A2(_03868_ ), .A3(_03822_ ), .A4(_03839_ ), .ZN(_03873_ ) );
OAI21_X1 _18059_ ( .A(\u_lsu.pmem[3297] ), .B1(_03864_ ), .B2(_10820_ ), .ZN(_03874_ ) );
AOI21_X1 _18060_ ( .A(fanout_net_48 ), .B1(_03873_ ), .B2(_03874_ ), .ZN(_01383_ ) );
BUF_X8 _18061_ ( .A(_09877_ ), .Z(_03875_ ) );
BUF_X4 _18062_ ( .A(_03875_ ), .Z(_03876_ ) );
NAND4_X1 _18063_ ( .A1(_09791_ ), .A2(_03868_ ), .A3(_03876_ ), .A4(_03839_ ), .ZN(_03877_ ) );
OAI21_X1 _18064_ ( .A(\u_lsu.pmem[3296] ), .B1(_03864_ ), .B2(_10820_ ), .ZN(_03878_ ) );
AOI21_X1 _18065_ ( .A(fanout_net_48 ), .B1(_03877_ ), .B2(_03878_ ), .ZN(_01384_ ) );
NAND4_X1 _18066_ ( .A1(_03793_ ), .A2(_02935_ ), .A3(_09914_ ), .A4(_10847_ ), .ZN(_03879_ ) );
OAI21_X1 _18067_ ( .A(\u_lsu.pmem[3271] ), .B1(_03864_ ), .B2(_10849_ ), .ZN(_03880_ ) );
AOI21_X1 _18068_ ( .A(fanout_net_48 ), .B1(_03879_ ), .B2(_03880_ ), .ZN(_01385_ ) );
NAND4_X1 _18069_ ( .A1(_09804_ ), .A2(_10974_ ), .A3(\alu_result_out[8] ), .A4(_10585_ ), .ZN(_03881_ ) );
OAI21_X1 _18070_ ( .A(\u_lsu.pmem[3270] ), .B1(_03864_ ), .B2(_10849_ ), .ZN(_03882_ ) );
AOI21_X1 _18071_ ( .A(fanout_net_48 ), .B1(_03881_ ), .B2(_03882_ ), .ZN(_01386_ ) );
NAND4_X1 _18072_ ( .A1(_09811_ ), .A2(_03735_ ), .A3(_03876_ ), .A4(_03839_ ), .ZN(_03883_ ) );
OAI21_X1 _18073_ ( .A(\u_lsu.pmem[3269] ), .B1(_03864_ ), .B2(_10848_ ), .ZN(_03884_ ) );
AOI21_X1 _18074_ ( .A(fanout_net_48 ), .B1(_03883_ ), .B2(_03884_ ), .ZN(_01387_ ) );
BUF_X4 _18075_ ( .A(_03396_ ), .Z(_03885_ ) );
BUF_X4 _18076_ ( .A(_03326_ ), .Z(_03886_ ) );
NAND4_X1 _18077_ ( .A1(_09835_ ), .A2(_03885_ ), .A3(_03886_ ), .A4(_03834_ ), .ZN(_03887_ ) );
OAI21_X1 _18078_ ( .A(\u_lsu.pmem[4288] ), .B1(_03810_ ), .B2(_09799_ ), .ZN(_03888_ ) );
AOI21_X1 _18079_ ( .A(fanout_net_48 ), .B1(_03887_ ), .B2(_03888_ ), .ZN(_01388_ ) );
BUF_X4 _18080_ ( .A(_11492_ ), .Z(_03889_ ) );
NAND4_X1 _18081_ ( .A1(_09815_ ), .A2(_03735_ ), .A3(_03876_ ), .A4(_03889_ ), .ZN(_03890_ ) );
OAI21_X1 _18082_ ( .A(\u_lsu.pmem[3268] ), .B1(_03864_ ), .B2(_10848_ ), .ZN(_03891_ ) );
AOI21_X1 _18083_ ( .A(fanout_net_48 ), .B1(_03890_ ), .B2(_03891_ ), .ZN(_01389_ ) );
NAND4_X1 _18084_ ( .A1(_09819_ ), .A2(_03735_ ), .A3(_03876_ ), .A4(_03889_ ), .ZN(_03892_ ) );
BUF_X4 _18085_ ( .A(_09562_ ), .Z(_03893_ ) );
OAI21_X1 _18086_ ( .A(\u_lsu.pmem[3267] ), .B1(_03893_ ), .B2(_10848_ ), .ZN(_03894_ ) );
AOI21_X1 _18087_ ( .A(fanout_net_48 ), .B1(_03892_ ), .B2(_03894_ ), .ZN(_01390_ ) );
NAND4_X1 _18088_ ( .A1(_09827_ ), .A2(_03868_ ), .A3(_03876_ ), .A4(_03889_ ), .ZN(_03895_ ) );
OAI21_X1 _18089_ ( .A(\u_lsu.pmem[3266] ), .B1(_03893_ ), .B2(_10848_ ), .ZN(_03896_ ) );
AOI21_X1 _18090_ ( .A(fanout_net_48 ), .B1(_03895_ ), .B2(_03896_ ), .ZN(_01391_ ) );
NAND4_X1 _18091_ ( .A1(_09831_ ), .A2(_03868_ ), .A3(_03876_ ), .A4(_03889_ ), .ZN(_03897_ ) );
OAI21_X1 _18092_ ( .A(\u_lsu.pmem[3265] ), .B1(_03893_ ), .B2(_10848_ ), .ZN(_03898_ ) );
AOI21_X1 _18093_ ( .A(fanout_net_48 ), .B1(_03897_ ), .B2(_03898_ ), .ZN(_01392_ ) );
NAND4_X1 _18094_ ( .A1(_09835_ ), .A2(_03868_ ), .A3(_03876_ ), .A4(_03889_ ), .ZN(_03899_ ) );
OAI21_X1 _18095_ ( .A(\u_lsu.pmem[3264] ), .B1(_03893_ ), .B2(_10848_ ), .ZN(_03900_ ) );
AOI21_X1 _18096_ ( .A(fanout_net_48 ), .B1(_03899_ ), .B2(_03900_ ), .ZN(_01393_ ) );
NAND4_X1 _18097_ ( .A1(_09840_ ), .A2(_03868_ ), .A3(_03876_ ), .A4(_03889_ ), .ZN(_03901_ ) );
OAI21_X1 _18098_ ( .A(\u_lsu.pmem[3239] ), .B1(_03893_ ), .B2(_10871_ ), .ZN(_03902_ ) );
AOI21_X1 _18099_ ( .A(fanout_net_49 ), .B1(_03901_ ), .B2(_03902_ ), .ZN(_01394_ ) );
NAND4_X1 _18100_ ( .A1(_09849_ ), .A2(_10974_ ), .A3(_10876_ ), .A4(_03674_ ), .ZN(_03903_ ) );
OAI21_X1 _18101_ ( .A(\u_lsu.pmem[3238] ), .B1(_03893_ ), .B2(_10871_ ), .ZN(_03904_ ) );
AOI21_X1 _18102_ ( .A(fanout_net_49 ), .B1(_03903_ ), .B2(_03904_ ), .ZN(_01395_ ) );
NAND4_X1 _18103_ ( .A1(_09853_ ), .A2(_03868_ ), .A3(_03876_ ), .A4(_03889_ ), .ZN(_03905_ ) );
OAI21_X1 _18104_ ( .A(\u_lsu.pmem[3237] ), .B1(_03893_ ), .B2(_10870_ ), .ZN(_03906_ ) );
AOI21_X1 _18105_ ( .A(fanout_net_49 ), .B1(_03905_ ), .B2(_03906_ ), .ZN(_01396_ ) );
NAND4_X1 _18106_ ( .A1(_09858_ ), .A2(_03868_ ), .A3(_03876_ ), .A4(_03889_ ), .ZN(_03907_ ) );
OAI21_X1 _18107_ ( .A(\u_lsu.pmem[3236] ), .B1(_03893_ ), .B2(_10870_ ), .ZN(_03908_ ) );
AOI21_X1 _18108_ ( .A(fanout_net_49 ), .B1(_03907_ ), .B2(_03908_ ), .ZN(_01397_ ) );
BUF_X4 _18109_ ( .A(_03020_ ), .Z(_03909_ ) );
BUF_X4 _18110_ ( .A(_03875_ ), .Z(_03910_ ) );
NAND4_X1 _18111_ ( .A1(_09861_ ), .A2(_03909_ ), .A3(_03910_ ), .A4(_03889_ ), .ZN(_03911_ ) );
OAI21_X1 _18112_ ( .A(\u_lsu.pmem[3235] ), .B1(_03893_ ), .B2(_10870_ ), .ZN(_03912_ ) );
AOI21_X1 _18113_ ( .A(fanout_net_49 ), .B1(_03911_ ), .B2(_03912_ ), .ZN(_01398_ ) );
NAND4_X1 _18114_ ( .A1(_09840_ ), .A2(_03885_ ), .A3(_03886_ ), .A4(_03834_ ), .ZN(_03913_ ) );
OAI21_X1 _18115_ ( .A(\u_lsu.pmem[4263] ), .B1(_03810_ ), .B2(_09846_ ), .ZN(_03914_ ) );
AOI21_X1 _18116_ ( .A(fanout_net_49 ), .B1(_03913_ ), .B2(_03914_ ), .ZN(_01399_ ) );
NAND4_X1 _18117_ ( .A1(_09864_ ), .A2(_03909_ ), .A3(_03910_ ), .A4(_03889_ ), .ZN(_03915_ ) );
OAI21_X1 _18118_ ( .A(\u_lsu.pmem[3234] ), .B1(_03893_ ), .B2(_10870_ ), .ZN(_03916_ ) );
AOI21_X1 _18119_ ( .A(fanout_net_49 ), .B1(_03915_ ), .B2(_03916_ ), .ZN(_01400_ ) );
BUF_X4 _18120_ ( .A(_11492_ ), .Z(_03917_ ) );
NAND4_X1 _18121_ ( .A1(_09867_ ), .A2(_03909_ ), .A3(_03910_ ), .A4(_03917_ ), .ZN(_03918_ ) );
BUF_X8 _18122_ ( .A(_09471_ ), .Z(_03919_ ) );
BUF_X4 _18123_ ( .A(_03919_ ), .Z(_03920_ ) );
OAI21_X1 _18124_ ( .A(\u_lsu.pmem[3233] ), .B1(_03920_ ), .B2(_10870_ ), .ZN(_03921_ ) );
AOI21_X1 _18125_ ( .A(fanout_net_49 ), .B1(_03918_ ), .B2(_03921_ ), .ZN(_01401_ ) );
NAND4_X1 _18126_ ( .A1(_09881_ ), .A2(_03735_ ), .A3(_03910_ ), .A4(_03917_ ), .ZN(_03922_ ) );
OAI21_X1 _18127_ ( .A(\u_lsu.pmem[3232] ), .B1(_03920_ ), .B2(_10870_ ), .ZN(_03923_ ) );
AOI21_X1 _18128_ ( .A(fanout_net_49 ), .B1(_03922_ ), .B2(_03923_ ), .ZN(_01402_ ) );
OAI21_X1 _18129_ ( .A(\u_lsu.pmem[3207] ), .B1(_10896_ ), .B2(_03769_ ), .ZN(_03924_ ) );
BUF_X4 _18130_ ( .A(_09522_ ), .Z(_03925_ ) );
NAND4_X1 _18131_ ( .A1(_03063_ ), .A2(_03478_ ), .A3(_02672_ ), .A4(_03925_ ), .ZN(_03926_ ) );
AOI21_X1 _18132_ ( .A(fanout_net_49 ), .B1(_03924_ ), .B2(_03926_ ), .ZN(_01403_ ) );
OAI21_X1 _18133_ ( .A(\u_lsu.pmem[3206] ), .B1(_10896_ ), .B2(_03769_ ), .ZN(_03927_ ) );
BUF_X4 _18134_ ( .A(_11381_ ), .Z(_03928_ ) );
NAND4_X1 _18135_ ( .A1(_03063_ ), .A2(_03056_ ), .A3(_03928_ ), .A4(_03925_ ), .ZN(_03929_ ) );
AOI21_X1 _18136_ ( .A(fanout_net_49 ), .B1(_03927_ ), .B2(_03929_ ), .ZN(_01404_ ) );
OAI21_X1 _18137_ ( .A(\u_lsu.pmem[3205] ), .B1(_10895_ ), .B2(_03769_ ), .ZN(_03930_ ) );
NAND4_X1 _18138_ ( .A1(_03063_ ), .A2(_03059_ ), .A3(_03928_ ), .A4(_03925_ ), .ZN(_03931_ ) );
AOI21_X1 _18139_ ( .A(fanout_net_49 ), .B1(_03930_ ), .B2(_03931_ ), .ZN(_01405_ ) );
BUF_X4 _18140_ ( .A(_09647_ ), .Z(_03932_ ) );
OAI21_X1 _18141_ ( .A(\u_lsu.pmem[3204] ), .B1(_10895_ ), .B2(_03932_ ), .ZN(_03933_ ) );
NAND4_X1 _18142_ ( .A1(_03063_ ), .A2(_03064_ ), .A3(_03928_ ), .A4(_03925_ ), .ZN(_03934_ ) );
AOI21_X1 _18143_ ( .A(fanout_net_49 ), .B1(_03933_ ), .B2(_03934_ ), .ZN(_01406_ ) );
OAI21_X1 _18144_ ( .A(\u_lsu.pmem[3203] ), .B1(_10895_ ), .B2(_03932_ ), .ZN(_03935_ ) );
NAND4_X1 _18145_ ( .A1(_03063_ ), .A2(_10915_ ), .A3(_03928_ ), .A4(_03925_ ), .ZN(_03936_ ) );
AOI21_X1 _18146_ ( .A(fanout_net_49 ), .B1(_03935_ ), .B2(_03936_ ), .ZN(_01407_ ) );
OAI21_X1 _18147_ ( .A(\u_lsu.pmem[3202] ), .B1(_10895_ ), .B2(_03932_ ), .ZN(_03937_ ) );
NAND4_X1 _18148_ ( .A1(_09906_ ), .A2(_03107_ ), .A3(_03928_ ), .A4(_03925_ ), .ZN(_03938_ ) );
AOI21_X1 _18149_ ( .A(fanout_net_49 ), .B1(_03937_ ), .B2(_03938_ ), .ZN(_01408_ ) );
OAI21_X1 _18150_ ( .A(\u_lsu.pmem[3201] ), .B1(_10895_ ), .B2(_03932_ ), .ZN(_03939_ ) );
NAND4_X1 _18151_ ( .A1(_03063_ ), .A2(_02308_ ), .A3(_03928_ ), .A4(_03925_ ), .ZN(_03940_ ) );
AOI21_X1 _18152_ ( .A(fanout_net_49 ), .B1(_03939_ ), .B2(_03940_ ), .ZN(_01409_ ) );
OAI21_X1 _18153_ ( .A(\u_lsu.pmem[4385] ), .B1(_09441_ ), .B2(_03666_ ), .ZN(_03941_ ) );
NAND4_X1 _18154_ ( .A1(_03143_ ), .A2(_03504_ ), .A3(_09131_ ), .A4(_09456_ ), .ZN(_03942_ ) );
AOI21_X1 _18155_ ( .A(fanout_net_49 ), .B1(_03941_ ), .B2(_03942_ ), .ZN(_01410_ ) );
NAND4_X1 _18156_ ( .A1(_09849_ ), .A2(_03885_ ), .A3(_03886_ ), .A4(_03834_ ), .ZN(_03943_ ) );
OAI21_X1 _18157_ ( .A(\u_lsu.pmem[4262] ), .B1(_03810_ ), .B2(_09846_ ), .ZN(_03944_ ) );
AOI21_X1 _18158_ ( .A(fanout_net_49 ), .B1(_03943_ ), .B2(_03944_ ), .ZN(_01411_ ) );
OAI21_X1 _18159_ ( .A(\u_lsu.pmem[3200] ), .B1(_10895_ ), .B2(_03932_ ), .ZN(_03945_ ) );
NAND4_X1 _18160_ ( .A1(_10898_ ), .A2(_11131_ ), .A3(_03928_ ), .A4(_03925_ ), .ZN(_03946_ ) );
AOI21_X1 _18161_ ( .A(fanout_net_49 ), .B1(_03945_ ), .B2(_03946_ ), .ZN(_01412_ ) );
AND2_X1 _18162_ ( .A1(_10925_ ), .A2(_10012_ ), .ZN(_03947_ ) );
OAI21_X1 _18163_ ( .A(_10715_ ), .B1(_03947_ ), .B2(\u_lsu.pmem[3175] ), .ZN(_03948_ ) );
AOI21_X1 _18164_ ( .A(_03948_ ), .B1(_09638_ ), .B2(_03947_ ), .ZN(_01413_ ) );
OAI21_X1 _18165_ ( .A(\u_lsu.pmem[3174] ), .B1(_10927_ ), .B2(\alu_result_out[9] ), .ZN(_03949_ ) );
BUF_X4 _18166_ ( .A(_09443_ ), .Z(_03950_ ) );
NAND4_X1 _18167_ ( .A1(_03950_ ), .A2(_09578_ ), .A3(_03928_ ), .A4(_10929_ ), .ZN(_03951_ ) );
AOI21_X1 _18168_ ( .A(fanout_net_49 ), .B1(_03949_ ), .B2(_03951_ ), .ZN(_01414_ ) );
OAI21_X1 _18169_ ( .A(\u_lsu.pmem[3173] ), .B1(_10927_ ), .B2(\alu_result_out[9] ), .ZN(_03952_ ) );
NAND4_X1 _18170_ ( .A1(_03950_ ), .A2(_09585_ ), .A3(_03928_ ), .A4(_10929_ ), .ZN(_03953_ ) );
AOI21_X1 _18171_ ( .A(fanout_net_49 ), .B1(_03952_ ), .B2(_03953_ ), .ZN(_01415_ ) );
OAI21_X1 _18172_ ( .A(\u_lsu.pmem[3172] ), .B1(_10926_ ), .B2(\alu_result_out[9] ), .ZN(_03954_ ) );
NAND4_X1 _18173_ ( .A1(_03950_ ), .A2(_11151_ ), .A3(_03928_ ), .A4(_10929_ ), .ZN(_03955_ ) );
AOI21_X1 _18174_ ( .A(fanout_net_49 ), .B1(_03954_ ), .B2(_03955_ ), .ZN(_01416_ ) );
OAI21_X1 _18175_ ( .A(\u_lsu.pmem[3171] ), .B1(_10926_ ), .B2(\alu_result_out[9] ), .ZN(_03956_ ) );
BUF_X4 _18176_ ( .A(_09443_ ), .Z(_03957_ ) );
BUF_X4 _18177_ ( .A(_11381_ ), .Z(_03958_ ) );
NAND4_X1 _18178_ ( .A1(_03957_ ), .A2(_09934_ ), .A3(_03958_ ), .A4(_10929_ ), .ZN(_03959_ ) );
AOI21_X1 _18179_ ( .A(fanout_net_49 ), .B1(_03956_ ), .B2(_03959_ ), .ZN(_01417_ ) );
OAI21_X1 _18180_ ( .A(\u_lsu.pmem[3170] ), .B1(_10926_ ), .B2(_10576_ ), .ZN(_03960_ ) );
NAND4_X1 _18181_ ( .A1(_03957_ ), .A2(_10015_ ), .A3(_03958_ ), .A4(_10929_ ), .ZN(_03961_ ) );
AOI21_X1 _18182_ ( .A(fanout_net_49 ), .B1(_03960_ ), .B2(_03961_ ), .ZN(_01418_ ) );
OAI21_X1 _18183_ ( .A(\u_lsu.pmem[3169] ), .B1(_10926_ ), .B2(_10576_ ), .ZN(_03962_ ) );
NAND4_X1 _18184_ ( .A1(_03957_ ), .A2(_09941_ ), .A3(_03958_ ), .A4(_10929_ ), .ZN(_03963_ ) );
AOI21_X1 _18185_ ( .A(fanout_net_49 ), .B1(_03962_ ), .B2(_03963_ ), .ZN(_01419_ ) );
OAI21_X1 _18186_ ( .A(\u_lsu.pmem[3168] ), .B1(_10926_ ), .B2(_10576_ ), .ZN(_03964_ ) );
NAND4_X1 _18187_ ( .A1(_03957_ ), .A2(_09621_ ), .A3(_03958_ ), .A4(_10929_ ), .ZN(_03965_ ) );
AOI21_X1 _18188_ ( .A(fanout_net_49 ), .B1(_03964_ ), .B2(_03965_ ), .ZN(_01420_ ) );
AND2_X1 _18189_ ( .A1(_10954_ ), .A2(_10012_ ), .ZN(_03966_ ) );
OAI21_X1 _18190_ ( .A(_09109_ ), .B1(_03966_ ), .B2(\u_lsu.pmem[3143] ), .ZN(_03967_ ) );
AOI21_X1 _18191_ ( .A(_03967_ ), .B1(_09638_ ), .B2(_03966_ ), .ZN(_01421_ ) );
NAND4_X1 _18192_ ( .A1(_09853_ ), .A2(_03885_ ), .A3(_03886_ ), .A4(_03834_ ), .ZN(_03968_ ) );
OAI21_X1 _18193_ ( .A(\u_lsu.pmem[4261] ), .B1(_03810_ ), .B2(_09845_ ), .ZN(_03969_ ) );
AOI21_X1 _18194_ ( .A(fanout_net_49 ), .B1(_03968_ ), .B2(_03969_ ), .ZN(_01422_ ) );
BUF_X4 _18195_ ( .A(_09953_ ), .Z(_03970_ ) );
NAND4_X1 _18196_ ( .A1(_03970_ ), .A2(_09957_ ), .A3(_03673_ ), .A4(_03674_ ), .ZN(_03971_ ) );
OAI21_X1 _18197_ ( .A(\u_lsu.pmem[3142] ), .B1(_10956_ ), .B2(_02584_ ), .ZN(_03972_ ) );
AOI21_X1 _18198_ ( .A(fanout_net_49 ), .B1(_03971_ ), .B2(_03972_ ), .ZN(_01423_ ) );
NAND4_X1 _18199_ ( .A1(_03970_ ), .A2(_09961_ ), .A3(_03673_ ), .A4(_03674_ ), .ZN(_03973_ ) );
BUF_X4 _18200_ ( .A(_09730_ ), .Z(_03974_ ) );
OAI21_X1 _18201_ ( .A(\u_lsu.pmem[3141] ), .B1(_10956_ ), .B2(_03974_ ), .ZN(_03975_ ) );
AOI21_X1 _18202_ ( .A(fanout_net_49 ), .B1(_03973_ ), .B2(_03975_ ), .ZN(_01424_ ) );
NAND4_X1 _18203_ ( .A1(_03970_ ), .A2(_09966_ ), .A3(_03673_ ), .A4(_03674_ ), .ZN(_03976_ ) );
OAI21_X1 _18204_ ( .A(\u_lsu.pmem[3140] ), .B1(_10955_ ), .B2(_03974_ ), .ZN(_03977_ ) );
AOI21_X1 _18205_ ( .A(fanout_net_49 ), .B1(_03976_ ), .B2(_03977_ ), .ZN(_01425_ ) );
BUF_X4 _18206_ ( .A(_10578_ ), .Z(_03978_ ) );
NAND4_X1 _18207_ ( .A1(_03970_ ), .A2(_09970_ ), .A3(_03673_ ), .A4(_03978_ ), .ZN(_03979_ ) );
OAI21_X1 _18208_ ( .A(\u_lsu.pmem[3139] ), .B1(_10955_ ), .B2(_03974_ ), .ZN(_03980_ ) );
AOI21_X1 _18209_ ( .A(fanout_net_50 ), .B1(_03979_ ), .B2(_03980_ ), .ZN(_01426_ ) );
NAND4_X1 _18210_ ( .A1(_03970_ ), .A2(_09974_ ), .A3(_03673_ ), .A4(_03978_ ), .ZN(_03981_ ) );
OAI21_X1 _18211_ ( .A(\u_lsu.pmem[3138] ), .B1(_10955_ ), .B2(_03974_ ), .ZN(_03982_ ) );
AOI21_X1 _18212_ ( .A(fanout_net_50 ), .B1(_03981_ ), .B2(_03982_ ), .ZN(_01427_ ) );
NAND4_X1 _18213_ ( .A1(_03970_ ), .A2(_09978_ ), .A3(_03673_ ), .A4(_03978_ ), .ZN(_03983_ ) );
OAI21_X1 _18214_ ( .A(\u_lsu.pmem[3137] ), .B1(_10955_ ), .B2(_03974_ ), .ZN(_03984_ ) );
AOI21_X1 _18215_ ( .A(fanout_net_50 ), .B1(_03983_ ), .B2(_03984_ ), .ZN(_01428_ ) );
NAND4_X1 _18216_ ( .A1(_03970_ ), .A2(_09982_ ), .A3(_03673_ ), .A4(_03978_ ), .ZN(_03985_ ) );
OAI21_X1 _18217_ ( .A(\u_lsu.pmem[3136] ), .B1(_10955_ ), .B2(_03974_ ), .ZN(_03986_ ) );
AOI21_X1 _18218_ ( .A(fanout_net_50 ), .B1(_03985_ ), .B2(_03986_ ), .ZN(_01429_ ) );
NAND4_X1 _18219_ ( .A1(_09987_ ), .A2(_03909_ ), .A3(_03910_ ), .A4(_03917_ ), .ZN(_03987_ ) );
NAND2_X1 _18220_ ( .A1(_09515_ ), .A2(_10980_ ), .ZN(_03988_ ) );
NAND2_X1 _18221_ ( .A1(_03988_ ), .A2(\u_lsu.pmem[3111] ), .ZN(_03989_ ) );
AOI21_X1 _18222_ ( .A(fanout_net_50 ), .B1(_03987_ ), .B2(_03989_ ), .ZN(_01430_ ) );
NAND4_X1 _18223_ ( .A1(_09994_ ), .A2(_03909_ ), .A3(_03910_ ), .A4(_03917_ ), .ZN(_03990_ ) );
NAND2_X1 _18224_ ( .A1(_03988_ ), .A2(\u_lsu.pmem[3110] ), .ZN(_03991_ ) );
AOI21_X1 _18225_ ( .A(fanout_net_50 ), .B1(_03990_ ), .B2(_03991_ ), .ZN(_01431_ ) );
NAND4_X1 _18226_ ( .A1(_09997_ ), .A2(_03909_ ), .A3(_03910_ ), .A4(_03917_ ), .ZN(_03992_ ) );
NAND2_X1 _18227_ ( .A1(_03988_ ), .A2(\u_lsu.pmem[3109] ), .ZN(_03993_ ) );
AOI21_X1 _18228_ ( .A(fanout_net_50 ), .B1(_03992_ ), .B2(_03993_ ), .ZN(_01432_ ) );
NAND4_X1 _18229_ ( .A1(_09858_ ), .A2(_03885_ ), .A3(_03886_ ), .A4(_03834_ ), .ZN(_03994_ ) );
OAI21_X1 _18230_ ( .A(\u_lsu.pmem[4260] ), .B1(_03810_ ), .B2(_09845_ ), .ZN(_03995_ ) );
AOI21_X1 _18231_ ( .A(fanout_net_50 ), .B1(_03994_ ), .B2(_03995_ ), .ZN(_01433_ ) );
NAND2_X1 _18232_ ( .A1(_03988_ ), .A2(\u_lsu.pmem[3108] ), .ZN(_03996_ ) );
NAND4_X1 _18233_ ( .A1(_03957_ ), .A2(_11151_ ), .A3(_03958_ ), .A4(_10979_ ), .ZN(_03997_ ) );
AOI21_X1 _18234_ ( .A(fanout_net_50 ), .B1(_03996_ ), .B2(_03997_ ), .ZN(_01434_ ) );
NAND2_X1 _18235_ ( .A1(_03988_ ), .A2(\u_lsu.pmem[3107] ), .ZN(_03998_ ) );
NAND4_X1 _18236_ ( .A1(_03957_ ), .A2(_09934_ ), .A3(_03958_ ), .A4(_10979_ ), .ZN(_03999_ ) );
AOI21_X1 _18237_ ( .A(fanout_net_50 ), .B1(_03998_ ), .B2(_03999_ ), .ZN(_01435_ ) );
NAND2_X1 _18238_ ( .A1(_03988_ ), .A2(\u_lsu.pmem[3106] ), .ZN(_04000_ ) );
NAND4_X1 _18239_ ( .A1(_03957_ ), .A2(_10015_ ), .A3(_03958_ ), .A4(_10979_ ), .ZN(_04001_ ) );
AOI21_X1 _18240_ ( .A(fanout_net_50 ), .B1(_04000_ ), .B2(_04001_ ), .ZN(_01436_ ) );
NAND2_X1 _18241_ ( .A1(_03988_ ), .A2(\u_lsu.pmem[3105] ), .ZN(_04002_ ) );
NAND4_X1 _18242_ ( .A1(_03957_ ), .A2(_09941_ ), .A3(_03958_ ), .A4(_10979_ ), .ZN(_04003_ ) );
AOI21_X1 _18243_ ( .A(fanout_net_50 ), .B1(_04002_ ), .B2(_04003_ ), .ZN(_01437_ ) );
NAND4_X1 _18244_ ( .A1(_10021_ ), .A2(_03909_ ), .A3(_03910_ ), .A4(_03917_ ), .ZN(_04004_ ) );
NAND2_X1 _18245_ ( .A1(_03988_ ), .A2(\u_lsu.pmem[3104] ), .ZN(_04005_ ) );
AOI21_X1 _18246_ ( .A(fanout_net_50 ), .B1(_04004_ ), .B2(_04005_ ), .ZN(_01438_ ) );
NAND4_X1 _18247_ ( .A1(_09700_ ), .A2(_11423_ ), .A3(_10974_ ), .A4(_11003_ ), .ZN(_04006_ ) );
OAI21_X1 _18248_ ( .A(\u_lsu.pmem[3079] ), .B1(_11006_ ), .B2(_03796_ ), .ZN(_04007_ ) );
AOI21_X1 _18249_ ( .A(fanout_net_50 ), .B1(_04006_ ), .B2(_04007_ ), .ZN(_01439_ ) );
BUF_X4 _18250_ ( .A(_09458_ ), .Z(_04008_ ) );
BUF_X4 _18251_ ( .A(_04008_ ), .Z(_04009_ ) );
NAND3_X1 _18252_ ( .A1(_04009_ ), .A2(_11145_ ), .A3(_11003_ ), .ZN(_04010_ ) );
OAI21_X1 _18253_ ( .A(\u_lsu.pmem[3078] ), .B1(_11006_ ), .B2(_03796_ ), .ZN(_04011_ ) );
AOI21_X1 _18254_ ( .A(fanout_net_50 ), .B1(_04010_ ), .B2(_04011_ ), .ZN(_01440_ ) );
NAND3_X1 _18255_ ( .A1(_04009_ ), .A2(_11148_ ), .A3(_11003_ ), .ZN(_04012_ ) );
BUF_X4 _18256_ ( .A(_10046_ ), .Z(_04013_ ) );
OAI21_X1 _18257_ ( .A(\u_lsu.pmem[3077] ), .B1(_11005_ ), .B2(_04013_ ), .ZN(_04014_ ) );
AOI21_X1 _18258_ ( .A(fanout_net_50 ), .B1(_04012_ ), .B2(_04014_ ), .ZN(_01441_ ) );
NAND3_X1 _18259_ ( .A1(_04009_ ), .A2(_03084_ ), .A3(_11003_ ), .ZN(_04015_ ) );
OAI21_X1 _18260_ ( .A(\u_lsu.pmem[3076] ), .B1(_11005_ ), .B2(_04013_ ), .ZN(_04016_ ) );
AOI21_X1 _18261_ ( .A(fanout_net_50 ), .B1(_04015_ ), .B2(_04016_ ), .ZN(_01442_ ) );
NAND3_X1 _18262_ ( .A1(_04009_ ), .A2(_03114_ ), .A3(_11003_ ), .ZN(_04017_ ) );
OAI21_X1 _18263_ ( .A(\u_lsu.pmem[3075] ), .B1(_11005_ ), .B2(_04013_ ), .ZN(_04018_ ) );
AOI21_X1 _18264_ ( .A(fanout_net_50 ), .B1(_04017_ ), .B2(_04018_ ), .ZN(_01443_ ) );
NAND4_X1 _18265_ ( .A1(_09861_ ), .A2(_03885_ ), .A3(_03886_ ), .A4(_03834_ ), .ZN(_04019_ ) );
OAI21_X1 _18266_ ( .A(\u_lsu.pmem[4259] ), .B1(_03810_ ), .B2(_09845_ ), .ZN(_04020_ ) );
AOI21_X1 _18267_ ( .A(fanout_net_50 ), .B1(_04019_ ), .B2(_04020_ ), .ZN(_01444_ ) );
NAND4_X1 _18268_ ( .A1(_11021_ ), .A2(_03885_ ), .A3(_03910_ ), .A4(_03917_ ), .ZN(_04021_ ) );
OAI21_X1 _18269_ ( .A(\u_lsu.pmem[3074] ), .B1(_11005_ ), .B2(_04013_ ), .ZN(_04022_ ) );
AOI21_X1 _18270_ ( .A(fanout_net_50 ), .B1(_04021_ ), .B2(_04022_ ), .ZN(_01445_ ) );
NAND3_X1 _18271_ ( .A1(_04009_ ), .A2(_03174_ ), .A3(_11003_ ), .ZN(_04023_ ) );
OAI21_X1 _18272_ ( .A(\u_lsu.pmem[3073] ), .B1(_11005_ ), .B2(_04013_ ), .ZN(_04024_ ) );
AOI21_X1 _18273_ ( .A(fanout_net_50 ), .B1(_04023_ ), .B2(_04024_ ), .ZN(_01446_ ) );
NAND3_X1 _18274_ ( .A1(_04009_ ), .A2(_03203_ ), .A3(_11003_ ), .ZN(_04025_ ) );
OAI21_X1 _18275_ ( .A(\u_lsu.pmem[3072] ), .B1(_11005_ ), .B2(_04013_ ), .ZN(_04026_ ) );
AOI21_X1 _18276_ ( .A(fanout_net_50 ), .B1(_04025_ ), .B2(_04026_ ), .ZN(_01447_ ) );
NOR2_X2 _18277_ ( .A1(_03850_ ), .A2(_11031_ ), .ZN(_04027_ ) );
NOR2_X1 _18278_ ( .A1(_04027_ ), .A2(\u_lsu.pmem[3047] ), .ZN(_04028_ ) );
AOI211_X1 _18279_ ( .A(fanout_net_50 ), .B(_04028_ ), .C1(_09568_ ), .C2(_04027_ ), .ZN(_01448_ ) );
NAND4_X1 _18280_ ( .A1(_10062_ ), .A2(_03885_ ), .A3(_03910_ ), .A4(_03917_ ), .ZN(_04029_ ) );
OAI21_X1 _18281_ ( .A(\u_lsu.pmem[3046] ), .B1(_03920_ ), .B2(_11032_ ), .ZN(_04030_ ) );
AOI21_X1 _18282_ ( .A(fanout_net_50 ), .B1(_04029_ ), .B2(_04030_ ), .ZN(_01449_ ) );
BUF_X4 _18283_ ( .A(_03875_ ), .Z(_04031_ ) );
NAND4_X1 _18284_ ( .A1(_10075_ ), .A2(_03885_ ), .A3(_04031_ ), .A4(_03917_ ), .ZN(_04032_ ) );
OAI21_X1 _18285_ ( .A(\u_lsu.pmem[3045] ), .B1(_03920_ ), .B2(_11032_ ), .ZN(_04033_ ) );
AOI21_X1 _18286_ ( .A(fanout_net_50 ), .B1(_04032_ ), .B2(_04033_ ), .ZN(_01450_ ) );
NAND4_X1 _18287_ ( .A1(_10079_ ), .A2(_03885_ ), .A3(_04031_ ), .A4(_03917_ ), .ZN(_04034_ ) );
OAI21_X1 _18288_ ( .A(\u_lsu.pmem[3044] ), .B1(_03920_ ), .B2(_11031_ ), .ZN(_04035_ ) );
AOI21_X1 _18289_ ( .A(fanout_net_50 ), .B1(_04034_ ), .B2(_04035_ ), .ZN(_01451_ ) );
BUF_X4 _18290_ ( .A(_03396_ ), .Z(_04036_ ) );
BUF_X4 _18291_ ( .A(_11492_ ), .Z(_04037_ ) );
NAND4_X1 _18292_ ( .A1(_10084_ ), .A2(_04036_ ), .A3(_04031_ ), .A4(_04037_ ), .ZN(_04038_ ) );
OAI21_X1 _18293_ ( .A(\u_lsu.pmem[3043] ), .B1(_03920_ ), .B2(_11031_ ), .ZN(_04039_ ) );
AOI21_X1 _18294_ ( .A(fanout_net_50 ), .B1(_04038_ ), .B2(_04039_ ), .ZN(_01452_ ) );
NAND4_X1 _18295_ ( .A1(_10088_ ), .A2(_04036_ ), .A3(_04031_ ), .A4(_04037_ ), .ZN(_04040_ ) );
OAI21_X1 _18296_ ( .A(\u_lsu.pmem[3042] ), .B1(_03920_ ), .B2(_11031_ ), .ZN(_04041_ ) );
AOI21_X1 _18297_ ( .A(fanout_net_50 ), .B1(_04040_ ), .B2(_04041_ ), .ZN(_01453_ ) );
NAND4_X1 _18298_ ( .A1(_10094_ ), .A2(_04036_ ), .A3(_04031_ ), .A4(_04037_ ), .ZN(_04042_ ) );
OAI21_X1 _18299_ ( .A(\u_lsu.pmem[3041] ), .B1(_03920_ ), .B2(_11031_ ), .ZN(_04043_ ) );
AOI21_X1 _18300_ ( .A(fanout_net_50 ), .B1(_04042_ ), .B2(_04043_ ), .ZN(_01454_ ) );
NAND4_X1 _18301_ ( .A1(_09864_ ), .A2(_04036_ ), .A3(_03886_ ), .A4(_03834_ ), .ZN(_04044_ ) );
OAI21_X1 _18302_ ( .A(\u_lsu.pmem[4258] ), .B1(_03810_ ), .B2(_09845_ ), .ZN(_04045_ ) );
AOI21_X1 _18303_ ( .A(fanout_net_50 ), .B1(_04044_ ), .B2(_04045_ ), .ZN(_01455_ ) );
NAND4_X1 _18304_ ( .A1(_10098_ ), .A2(_04036_ ), .A3(_04031_ ), .A4(_04037_ ), .ZN(_04046_ ) );
OAI21_X1 _18305_ ( .A(\u_lsu.pmem[3040] ), .B1(_03920_ ), .B2(_11031_ ), .ZN(_04047_ ) );
AOI21_X1 _18306_ ( .A(fanout_net_51 ), .B1(_04046_ ), .B2(_04047_ ), .ZN(_01456_ ) );
NOR2_X2 _18307_ ( .A1(_03850_ ), .A2(_11058_ ), .ZN(_04048_ ) );
NOR2_X1 _18308_ ( .A1(_04048_ ), .A2(\u_lsu.pmem[3015] ), .ZN(_04049_ ) );
AOI211_X1 _18309_ ( .A(fanout_net_51 ), .B(_04049_ ), .C1(_09568_ ), .C2(_04048_ ), .ZN(_01457_ ) );
NAND4_X1 _18310_ ( .A1(_10117_ ), .A2(_04036_ ), .A3(_04031_ ), .A4(_04037_ ), .ZN(_04050_ ) );
OAI21_X1 _18311_ ( .A(\u_lsu.pmem[3014] ), .B1(_03920_ ), .B2(_11059_ ), .ZN(_04051_ ) );
AOI21_X1 _18312_ ( .A(fanout_net_51 ), .B1(_04050_ ), .B2(_04051_ ), .ZN(_01458_ ) );
NAND4_X1 _18313_ ( .A1(_10121_ ), .A2(_04036_ ), .A3(_04031_ ), .A4(_04037_ ), .ZN(_04052_ ) );
BUF_X4 _18314_ ( .A(_03919_ ), .Z(_04053_ ) );
OAI21_X1 _18315_ ( .A(\u_lsu.pmem[3013] ), .B1(_04053_ ), .B2(_11059_ ), .ZN(_04054_ ) );
AOI21_X1 _18316_ ( .A(fanout_net_51 ), .B1(_04052_ ), .B2(_04054_ ), .ZN(_01459_ ) );
NAND4_X1 _18317_ ( .A1(_10125_ ), .A2(_04036_ ), .A3(_04031_ ), .A4(_04037_ ), .ZN(_04055_ ) );
OAI21_X1 _18318_ ( .A(\u_lsu.pmem[3012] ), .B1(_04053_ ), .B2(_11058_ ), .ZN(_04056_ ) );
AOI21_X1 _18319_ ( .A(fanout_net_51 ), .B1(_04055_ ), .B2(_04056_ ), .ZN(_01460_ ) );
NAND4_X1 _18320_ ( .A1(_10131_ ), .A2(_04036_ ), .A3(_04031_ ), .A4(_04037_ ), .ZN(_04057_ ) );
OAI21_X1 _18321_ ( .A(\u_lsu.pmem[3011] ), .B1(_04053_ ), .B2(_11058_ ), .ZN(_04058_ ) );
AOI21_X1 _18322_ ( .A(fanout_net_51 ), .B1(_04057_ ), .B2(_04058_ ), .ZN(_01461_ ) );
BUF_X4 _18323_ ( .A(_03875_ ), .Z(_04059_ ) );
NAND4_X1 _18324_ ( .A1(_10135_ ), .A2(_04036_ ), .A3(_04059_ ), .A4(_04037_ ), .ZN(_04060_ ) );
OAI21_X1 _18325_ ( .A(\u_lsu.pmem[3010] ), .B1(_04053_ ), .B2(_11058_ ), .ZN(_04061_ ) );
AOI21_X1 _18326_ ( .A(fanout_net_51 ), .B1(_04060_ ), .B2(_04061_ ), .ZN(_01462_ ) );
BUF_X4 _18327_ ( .A(_03396_ ), .Z(_04062_ ) );
NAND4_X1 _18328_ ( .A1(_10138_ ), .A2(_04062_ ), .A3(_04059_ ), .A4(_04037_ ), .ZN(_04063_ ) );
OAI21_X1 _18329_ ( .A(\u_lsu.pmem[3009] ), .B1(_04053_ ), .B2(_11058_ ), .ZN(_04064_ ) );
AOI21_X1 _18330_ ( .A(fanout_net_51 ), .B1(_04063_ ), .B2(_04064_ ), .ZN(_01463_ ) );
BUF_X4 _18331_ ( .A(_11492_ ), .Z(_04065_ ) );
NAND4_X1 _18332_ ( .A1(_10144_ ), .A2(_04062_ ), .A3(_04059_ ), .A4(_04065_ ), .ZN(_04066_ ) );
OAI21_X1 _18333_ ( .A(\u_lsu.pmem[3008] ), .B1(_04053_ ), .B2(_11058_ ), .ZN(_04067_ ) );
AOI21_X1 _18334_ ( .A(fanout_net_51 ), .B1(_04066_ ), .B2(_04067_ ), .ZN(_01464_ ) );
NAND4_X1 _18335_ ( .A1(_10148_ ), .A2(_04062_ ), .A3(_04059_ ), .A4(_04065_ ), .ZN(_04068_ ) );
OAI21_X1 _18336_ ( .A(\u_lsu.pmem[2983] ), .B1(_04053_ ), .B2(_11088_ ), .ZN(_04069_ ) );
AOI21_X1 _18337_ ( .A(fanout_net_51 ), .B1(_04068_ ), .B2(_04069_ ), .ZN(_01465_ ) );
NAND4_X1 _18338_ ( .A1(_09867_ ), .A2(_04062_ ), .A3(_03886_ ), .A4(_03834_ ), .ZN(_04070_ ) );
BUF_X4 _18339_ ( .A(_09443_ ), .Z(_04071_ ) );
OAI21_X1 _18340_ ( .A(\u_lsu.pmem[4257] ), .B1(_04071_ ), .B2(_09845_ ), .ZN(_04072_ ) );
AOI21_X1 _18341_ ( .A(fanout_net_51 ), .B1(_04070_ ), .B2(_04072_ ), .ZN(_01466_ ) );
NAND4_X1 _18342_ ( .A1(_10156_ ), .A2(_04062_ ), .A3(_04059_ ), .A4(_04065_ ), .ZN(_04073_ ) );
OAI21_X1 _18343_ ( .A(\u_lsu.pmem[2982] ), .B1(_04053_ ), .B2(_11088_ ), .ZN(_04074_ ) );
AOI21_X1 _18344_ ( .A(fanout_net_51 ), .B1(_04073_ ), .B2(_04074_ ), .ZN(_01467_ ) );
NAND4_X1 _18345_ ( .A1(_10160_ ), .A2(_04062_ ), .A3(_04059_ ), .A4(_04065_ ), .ZN(_04075_ ) );
OAI21_X1 _18346_ ( .A(\u_lsu.pmem[2981] ), .B1(_04053_ ), .B2(_11087_ ), .ZN(_04076_ ) );
AOI21_X1 _18347_ ( .A(fanout_net_51 ), .B1(_04075_ ), .B2(_04076_ ), .ZN(_01468_ ) );
NAND4_X1 _18348_ ( .A1(_10166_ ), .A2(_04062_ ), .A3(_04059_ ), .A4(_04065_ ), .ZN(_04077_ ) );
OAI21_X1 _18349_ ( .A(\u_lsu.pmem[2980] ), .B1(_04053_ ), .B2(_11087_ ), .ZN(_04078_ ) );
AOI21_X1 _18350_ ( .A(fanout_net_51 ), .B1(_04077_ ), .B2(_04078_ ), .ZN(_01469_ ) );
NAND4_X1 _18351_ ( .A1(_10169_ ), .A2(_04062_ ), .A3(_04059_ ), .A4(_04065_ ), .ZN(_04079_ ) );
BUF_X4 _18352_ ( .A(_03919_ ), .Z(_04080_ ) );
OAI21_X1 _18353_ ( .A(\u_lsu.pmem[2979] ), .B1(_04080_ ), .B2(_11087_ ), .ZN(_04081_ ) );
AOI21_X1 _18354_ ( .A(fanout_net_51 ), .B1(_04079_ ), .B2(_04081_ ), .ZN(_01470_ ) );
NAND4_X1 _18355_ ( .A1(_10172_ ), .A2(_04062_ ), .A3(_04059_ ), .A4(_04065_ ), .ZN(_04082_ ) );
OAI21_X1 _18356_ ( .A(\u_lsu.pmem[2978] ), .B1(_04080_ ), .B2(_11087_ ), .ZN(_04083_ ) );
AOI21_X1 _18357_ ( .A(fanout_net_51 ), .B1(_04082_ ), .B2(_04083_ ), .ZN(_01471_ ) );
NAND4_X1 _18358_ ( .A1(_10176_ ), .A2(_04062_ ), .A3(_04059_ ), .A4(_04065_ ), .ZN(_04084_ ) );
OAI21_X1 _18359_ ( .A(\u_lsu.pmem[2977] ), .B1(_04080_ ), .B2(_11087_ ), .ZN(_04085_ ) );
AOI21_X1 _18360_ ( .A(fanout_net_51 ), .B1(_04084_ ), .B2(_04085_ ), .ZN(_01472_ ) );
NAND4_X1 _18361_ ( .A1(_03970_ ), .A2(_02935_ ), .A3(_03753_ ), .A4(_11086_ ), .ZN(_04086_ ) );
OAI21_X1 _18362_ ( .A(\u_lsu.pmem[2976] ), .B1(_04080_ ), .B2(_11087_ ), .ZN(_04087_ ) );
AOI21_X1 _18363_ ( .A(fanout_net_51 ), .B1(_04086_ ), .B2(_04087_ ), .ZN(_01473_ ) );
OAI21_X1 _18364_ ( .A(\u_lsu.pmem[2951] ), .B1(_11110_ ), .B2(_03932_ ), .ZN(_04088_ ) );
NAND4_X1 _18365_ ( .A1(_03254_ ), .A2(_03478_ ), .A3(_03958_ ), .A4(_03925_ ), .ZN(_04089_ ) );
AOI21_X1 _18366_ ( .A(fanout_net_51 ), .B1(_04088_ ), .B2(_04089_ ), .ZN(_01474_ ) );
OAI21_X1 _18367_ ( .A(\u_lsu.pmem[2950] ), .B1(_11110_ ), .B2(_03932_ ), .ZN(_04090_ ) );
NAND4_X1 _18368_ ( .A1(_03254_ ), .A2(_03056_ ), .A3(_03958_ ), .A4(_03925_ ), .ZN(_04091_ ) );
AOI21_X1 _18369_ ( .A(fanout_net_51 ), .B1(_04090_ ), .B2(_04091_ ), .ZN(_01475_ ) );
OAI21_X1 _18370_ ( .A(\u_lsu.pmem[2949] ), .B1(_11109_ ), .B2(_03932_ ), .ZN(_04092_ ) );
BUF_X4 _18371_ ( .A(_11381_ ), .Z(_04093_ ) );
BUF_X4 _18372_ ( .A(_09522_ ), .Z(_04094_ ) );
NAND4_X1 _18373_ ( .A1(_03254_ ), .A2(_03059_ ), .A3(_04093_ ), .A4(_04094_ ), .ZN(_04095_ ) );
AOI21_X1 _18374_ ( .A(fanout_net_51 ), .B1(_04092_ ), .B2(_04095_ ), .ZN(_01476_ ) );
BUF_X4 _18375_ ( .A(_03396_ ), .Z(_04096_ ) );
BUF_X4 _18376_ ( .A(_09730_ ), .Z(_04097_ ) );
NAND4_X1 _18377_ ( .A1(_09881_ ), .A2(_04096_ ), .A3(_03886_ ), .A4(_04097_ ), .ZN(_04098_ ) );
OAI21_X1 _18378_ ( .A(\u_lsu.pmem[4256] ), .B1(_04071_ ), .B2(_09845_ ), .ZN(_04099_ ) );
AOI21_X1 _18379_ ( .A(fanout_net_51 ), .B1(_04098_ ), .B2(_04099_ ), .ZN(_01477_ ) );
OAI21_X1 _18380_ ( .A(\u_lsu.pmem[2948] ), .B1(_11109_ ), .B2(_03932_ ), .ZN(_04100_ ) );
NAND4_X1 _18381_ ( .A1(_03254_ ), .A2(_03064_ ), .A3(_04093_ ), .A4(_04094_ ), .ZN(_04101_ ) );
AOI21_X1 _18382_ ( .A(fanout_net_51 ), .B1(_04100_ ), .B2(_04101_ ), .ZN(_01478_ ) );
OAI21_X1 _18383_ ( .A(\u_lsu.pmem[2947] ), .B1(_11109_ ), .B2(_03932_ ), .ZN(_04102_ ) );
NAND4_X1 _18384_ ( .A1(_03254_ ), .A2(_09519_ ), .A3(_04093_ ), .A4(_04094_ ), .ZN(_04103_ ) );
AOI21_X1 _18385_ ( .A(fanout_net_51 ), .B1(_04102_ ), .B2(_04103_ ), .ZN(_01479_ ) );
BUF_X4 _18386_ ( .A(_09647_ ), .Z(_04104_ ) );
OAI21_X1 _18387_ ( .A(\u_lsu.pmem[2946] ), .B1(_11109_ ), .B2(_04104_ ), .ZN(_04105_ ) );
NAND4_X1 _18388_ ( .A1(_09874_ ), .A2(_03361_ ), .A3(_04093_ ), .A4(_04094_ ), .ZN(_04106_ ) );
AOI21_X1 _18389_ ( .A(fanout_net_51 ), .B1(_04105_ ), .B2(_04106_ ), .ZN(_01480_ ) );
OAI21_X1 _18390_ ( .A(\u_lsu.pmem[2945] ), .B1(_11109_ ), .B2(_04104_ ), .ZN(_04107_ ) );
NAND4_X1 _18391_ ( .A1(_03254_ ), .A2(_02308_ ), .A3(_04093_ ), .A4(_04094_ ), .ZN(_04108_ ) );
AOI21_X1 _18392_ ( .A(fanout_net_51 ), .B1(_04107_ ), .B2(_04108_ ), .ZN(_01481_ ) );
OAI21_X1 _18393_ ( .A(\u_lsu.pmem[2944] ), .B1(_11109_ ), .B2(_04104_ ), .ZN(_04109_ ) );
NAND4_X1 _18394_ ( .A1(_11112_ ), .A2(_11131_ ), .A3(_04093_ ), .A4(_04094_ ), .ZN(_04110_ ) );
AOI21_X1 _18395_ ( .A(fanout_net_51 ), .B1(_04109_ ), .B2(_04110_ ), .ZN(_01482_ ) );
OAI21_X1 _18396_ ( .A(\u_lsu.pmem[2919] ), .B1(_11136_ ), .B2(_04104_ ), .ZN(_04111_ ) );
NAND3_X1 _18397_ ( .A1(_03826_ ), .A2(_11000_ ), .A3(_11140_ ), .ZN(_04112_ ) );
AOI21_X1 _18398_ ( .A(fanout_net_51 ), .B1(_04111_ ), .B2(_04112_ ), .ZN(_01483_ ) );
OAI21_X1 _18399_ ( .A(\u_lsu.pmem[2918] ), .B1(_11136_ ), .B2(_04104_ ), .ZN(_04113_ ) );
NAND3_X1 _18400_ ( .A1(_03826_ ), .A2(_09579_ ), .A3(_11140_ ), .ZN(_04114_ ) );
AOI21_X1 _18401_ ( .A(fanout_net_51 ), .B1(_04113_ ), .B2(_04114_ ), .ZN(_01484_ ) );
OAI21_X1 _18402_ ( .A(\u_lsu.pmem[2917] ), .B1(_11136_ ), .B2(_04104_ ), .ZN(_04115_ ) );
NAND3_X1 _18403_ ( .A1(_03826_ ), .A2(_09586_ ), .A3(_11134_ ), .ZN(_04116_ ) );
AOI21_X1 _18404_ ( .A(fanout_net_51 ), .B1(_04115_ ), .B2(_04116_ ), .ZN(_01485_ ) );
OAI21_X1 _18405_ ( .A(\u_lsu.pmem[2916] ), .B1(_11136_ ), .B2(_04104_ ), .ZN(_04117_ ) );
NAND3_X1 _18406_ ( .A1(_03826_ ), .A2(_09589_ ), .A3(_11134_ ), .ZN(_04118_ ) );
AOI21_X1 _18407_ ( .A(fanout_net_52 ), .B1(_04117_ ), .B2(_04118_ ), .ZN(_01486_ ) );
OAI21_X1 _18408_ ( .A(\u_lsu.pmem[2915] ), .B1(_11136_ ), .B2(_04104_ ), .ZN(_04119_ ) );
NAND3_X1 _18409_ ( .A1(_03826_ ), .A2(_09592_ ), .A3(_11134_ ), .ZN(_04120_ ) );
AOI21_X1 _18410_ ( .A(fanout_net_52 ), .B1(_04119_ ), .B2(_04120_ ), .ZN(_01487_ ) );
OAI21_X1 _18411_ ( .A(\u_lsu.pmem[4231] ), .B1(_09891_ ), .B2(_03666_ ), .ZN(_04121_ ) );
NAND4_X1 _18412_ ( .A1(_02301_ ), .A2(_03478_ ), .A3(_03640_ ), .A4(_03646_ ), .ZN(_04122_ ) );
AOI21_X1 _18413_ ( .A(fanout_net_52 ), .B1(_04121_ ), .B2(_04122_ ), .ZN(_01488_ ) );
OAI21_X1 _18414_ ( .A(\u_lsu.pmem[2914] ), .B1(_11136_ ), .B2(_04104_ ), .ZN(_04123_ ) );
NAND3_X1 _18415_ ( .A1(_03826_ ), .A2(_09695_ ), .A3(_11134_ ), .ZN(_04124_ ) );
AOI21_X1 _18416_ ( .A(fanout_net_52 ), .B1(_04123_ ), .B2(_04124_ ), .ZN(_01489_ ) );
OAI21_X1 _18417_ ( .A(\u_lsu.pmem[2913] ), .B1(_11136_ ), .B2(_04104_ ), .ZN(_04125_ ) );
BUF_X4 _18418_ ( .A(_09641_ ), .Z(_04126_ ) );
NAND3_X1 _18419_ ( .A1(_04126_ ), .A2(_09617_ ), .A3(_11134_ ), .ZN(_04127_ ) );
AOI21_X1 _18420_ ( .A(fanout_net_52 ), .B1(_04125_ ), .B2(_04127_ ), .ZN(_01490_ ) );
BUF_X4 _18421_ ( .A(_09647_ ), .Z(_04128_ ) );
OAI21_X1 _18422_ ( .A(\u_lsu.pmem[2912] ), .B1(_11136_ ), .B2(_04128_ ), .ZN(_04129_ ) );
NAND3_X1 _18423_ ( .A1(_04126_ ), .A2(_09622_ ), .A3(_11134_ ), .ZN(_04130_ ) );
AOI21_X1 _18424_ ( .A(fanout_net_52 ), .B1(_04129_ ), .B2(_04130_ ), .ZN(_01491_ ) );
OAI21_X1 _18425_ ( .A(\u_lsu.pmem[2887] ), .B1(_11171_ ), .B2(_04128_ ), .ZN(_04131_ ) );
NAND3_X1 _18426_ ( .A1(_04126_ ), .A2(_11000_ ), .A3(_11173_ ), .ZN(_04132_ ) );
AOI21_X1 _18427_ ( .A(fanout_net_52 ), .B1(_04131_ ), .B2(_04132_ ), .ZN(_01492_ ) );
OAI21_X1 _18428_ ( .A(\u_lsu.pmem[2886] ), .B1(_11171_ ), .B2(_04128_ ), .ZN(_04133_ ) );
NAND3_X1 _18429_ ( .A1(_04126_ ), .A2(_09579_ ), .A3(_11173_ ), .ZN(_04134_ ) );
AOI21_X1 _18430_ ( .A(fanout_net_52 ), .B1(_04133_ ), .B2(_04134_ ), .ZN(_01493_ ) );
OAI21_X1 _18431_ ( .A(\u_lsu.pmem[2885] ), .B1(_11171_ ), .B2(_04128_ ), .ZN(_04135_ ) );
NAND3_X1 _18432_ ( .A1(_04126_ ), .A2(_09586_ ), .A3(_11169_ ), .ZN(_04136_ ) );
AOI21_X1 _18433_ ( .A(fanout_net_52 ), .B1(_04135_ ), .B2(_04136_ ), .ZN(_01494_ ) );
OAI21_X1 _18434_ ( .A(\u_lsu.pmem[2884] ), .B1(_11171_ ), .B2(_04128_ ), .ZN(_04137_ ) );
NAND3_X1 _18435_ ( .A1(_04126_ ), .A2(_09589_ ), .A3(_11169_ ), .ZN(_04138_ ) );
AOI21_X1 _18436_ ( .A(fanout_net_52 ), .B1(_04137_ ), .B2(_04138_ ), .ZN(_01495_ ) );
OAI21_X1 _18437_ ( .A(\u_lsu.pmem[2883] ), .B1(_11171_ ), .B2(_04128_ ), .ZN(_04139_ ) );
NAND3_X1 _18438_ ( .A1(_04126_ ), .A2(_09592_ ), .A3(_11169_ ), .ZN(_04140_ ) );
AOI21_X1 _18439_ ( .A(fanout_net_52 ), .B1(_04139_ ), .B2(_04140_ ), .ZN(_01496_ ) );
OAI21_X1 _18440_ ( .A(\u_lsu.pmem[2882] ), .B1(_11171_ ), .B2(_04128_ ), .ZN(_04141_ ) );
NAND3_X1 _18441_ ( .A1(_04126_ ), .A2(_09695_ ), .A3(_11169_ ), .ZN(_04142_ ) );
AOI21_X1 _18442_ ( .A(fanout_net_52 ), .B1(_04141_ ), .B2(_04142_ ), .ZN(_01497_ ) );
OAI21_X1 _18443_ ( .A(\u_lsu.pmem[2881] ), .B1(_11171_ ), .B2(_04128_ ), .ZN(_04143_ ) );
NAND3_X1 _18444_ ( .A1(_04126_ ), .A2(_09617_ ), .A3(_11169_ ), .ZN(_04144_ ) );
AOI21_X1 _18445_ ( .A(fanout_net_52 ), .B1(_04143_ ), .B2(_04144_ ), .ZN(_01498_ ) );
OAI21_X1 _18446_ ( .A(\u_lsu.pmem[4230] ), .B1(_09891_ ), .B2(_09882_ ), .ZN(_04145_ ) );
NAND4_X1 _18447_ ( .A1(_02301_ ), .A2(_03056_ ), .A3(_03640_ ), .A4(_03646_ ), .ZN(_04146_ ) );
AOI21_X1 _18448_ ( .A(fanout_net_52 ), .B1(_04145_ ), .B2(_04146_ ), .ZN(_01499_ ) );
OAI21_X1 _18449_ ( .A(\u_lsu.pmem[2880] ), .B1(_11171_ ), .B2(_04128_ ), .ZN(_04147_ ) );
NAND3_X1 _18450_ ( .A1(_04126_ ), .A2(_09622_ ), .A3(_11169_ ), .ZN(_04148_ ) );
AOI21_X1 _18451_ ( .A(fanout_net_52 ), .B1(_04147_ ), .B2(_04148_ ), .ZN(_01500_ ) );
BUF_X4 _18452_ ( .A(_03875_ ), .Z(_04149_ ) );
NAND4_X1 _18453_ ( .A1(_10250_ ), .A2(_04096_ ), .A3(_04149_ ), .A4(_04065_ ), .ZN(_04150_ ) );
OAI21_X1 _18454_ ( .A(\u_lsu.pmem[2855] ), .B1(_11209_ ), .B2(_03974_ ), .ZN(_04151_ ) );
AOI21_X1 _18455_ ( .A(fanout_net_52 ), .B1(_04150_ ), .B2(_04151_ ), .ZN(_01501_ ) );
NAND4_X1 _18456_ ( .A1(_10263_ ), .A2(_04096_ ), .A3(_04149_ ), .A4(_04065_ ), .ZN(_04152_ ) );
OAI21_X1 _18457_ ( .A(\u_lsu.pmem[2854] ), .B1(_11209_ ), .B2(_03974_ ), .ZN(_04153_ ) );
AOI21_X1 _18458_ ( .A(fanout_net_52 ), .B1(_04152_ ), .B2(_04153_ ), .ZN(_01502_ ) );
BUF_X8 _18459_ ( .A(_09442_ ), .Z(_04154_ ) );
BUF_X4 _18460_ ( .A(_04154_ ), .Z(_04155_ ) );
NAND4_X1 _18461_ ( .A1(_10267_ ), .A2(_04096_ ), .A3(_04149_ ), .A4(_04155_ ), .ZN(_04156_ ) );
OAI21_X1 _18462_ ( .A(\u_lsu.pmem[2853] ), .B1(_11209_ ), .B2(_03974_ ), .ZN(_04157_ ) );
AOI21_X1 _18463_ ( .A(fanout_net_52 ), .B1(_04156_ ), .B2(_04157_ ), .ZN(_01503_ ) );
NOR2_X1 _18464_ ( .A1(_11199_ ), .A2(_09635_ ), .ZN(_04158_ ) );
OAI21_X1 _18465_ ( .A(_09109_ ), .B1(_04158_ ), .B2(\u_lsu.pmem[2852] ), .ZN(_04159_ ) );
AOI21_X1 _18466_ ( .A(_04159_ ), .B1(_09691_ ), .B2(_04158_ ), .ZN(_01504_ ) );
OAI21_X1 _18467_ ( .A(\u_lsu.pmem[2851] ), .B1(_11209_ ), .B2(_04128_ ), .ZN(_04160_ ) );
BUF_X4 _18468_ ( .A(_09641_ ), .Z(_04161_ ) );
NAND3_X1 _18469_ ( .A1(_04161_ ), .A2(_09592_ ), .A3(_11198_ ), .ZN(_04162_ ) );
AOI21_X1 _18470_ ( .A(fanout_net_52 ), .B1(_04160_ ), .B2(_04162_ ), .ZN(_01505_ ) );
BUF_X4 _18471_ ( .A(_09647_ ), .Z(_04163_ ) );
OAI21_X1 _18472_ ( .A(\u_lsu.pmem[2850] ), .B1(_11209_ ), .B2(_04163_ ), .ZN(_04164_ ) );
NAND3_X1 _18473_ ( .A1(_04161_ ), .A2(_09695_ ), .A3(_11198_ ), .ZN(_04165_ ) );
AOI21_X1 _18474_ ( .A(fanout_net_52 ), .B1(_04164_ ), .B2(_04165_ ), .ZN(_01506_ ) );
OAI21_X1 _18475_ ( .A(\u_lsu.pmem[2849] ), .B1(_11209_ ), .B2(_04163_ ), .ZN(_04166_ ) );
NAND3_X1 _18476_ ( .A1(_04161_ ), .A2(_09617_ ), .A3(_11198_ ), .ZN(_04167_ ) );
AOI21_X1 _18477_ ( .A(fanout_net_52 ), .B1(_04166_ ), .B2(_04167_ ), .ZN(_01507_ ) );
NAND4_X1 _18478_ ( .A1(_10279_ ), .A2(_04096_ ), .A3(_04149_ ), .A4(_04155_ ), .ZN(_04168_ ) );
OAI21_X1 _18479_ ( .A(\u_lsu.pmem[2848] ), .B1(_11209_ ), .B2(_03974_ ), .ZN(_04169_ ) );
AOI21_X1 _18480_ ( .A(fanout_net_52 ), .B1(_04168_ ), .B2(_04169_ ), .ZN(_01508_ ) );
NAND4_X1 _18481_ ( .A1(_10285_ ), .A2(_04096_ ), .A3(_04149_ ), .A4(_04155_ ), .ZN(_04170_ ) );
OAI21_X1 _18482_ ( .A(\u_lsu.pmem[2823] ), .B1(_04080_ ), .B2(_11225_ ), .ZN(_04171_ ) );
AOI21_X1 _18483_ ( .A(fanout_net_52 ), .B1(_04170_ ), .B2(_04171_ ), .ZN(_01509_ ) );
OAI21_X1 _18484_ ( .A(\u_lsu.pmem[4229] ), .B1(_09890_ ), .B2(_09882_ ), .ZN(_04172_ ) );
NAND4_X1 _18485_ ( .A1(_02301_ ), .A2(_03059_ ), .A3(_03640_ ), .A4(_03646_ ), .ZN(_04173_ ) );
AOI21_X1 _18486_ ( .A(fanout_net_52 ), .B1(_04172_ ), .B2(_04173_ ), .ZN(_01510_ ) );
NAND4_X1 _18487_ ( .A1(_10295_ ), .A2(_04096_ ), .A3(_04149_ ), .A4(_04155_ ), .ZN(_04174_ ) );
OAI21_X1 _18488_ ( .A(\u_lsu.pmem[2822] ), .B1(_04080_ ), .B2(_11225_ ), .ZN(_04175_ ) );
AOI21_X1 _18489_ ( .A(fanout_net_52 ), .B1(_04174_ ), .B2(_04175_ ), .ZN(_01511_ ) );
NAND4_X1 _18490_ ( .A1(_10299_ ), .A2(_04096_ ), .A3(_04149_ ), .A4(_04155_ ), .ZN(_04176_ ) );
OAI21_X1 _18491_ ( .A(\u_lsu.pmem[2821] ), .B1(_04080_ ), .B2(_11224_ ), .ZN(_04177_ ) );
AOI21_X1 _18492_ ( .A(fanout_net_52 ), .B1(_04176_ ), .B2(_04177_ ), .ZN(_01512_ ) );
NAND4_X1 _18493_ ( .A1(_10306_ ), .A2(_04096_ ), .A3(_04149_ ), .A4(_04155_ ), .ZN(_04178_ ) );
OAI21_X1 _18494_ ( .A(\u_lsu.pmem[2820] ), .B1(_04080_ ), .B2(_11224_ ), .ZN(_04179_ ) );
AOI21_X1 _18495_ ( .A(fanout_net_52 ), .B1(_04178_ ), .B2(_04179_ ), .ZN(_01513_ ) );
NAND4_X1 _18496_ ( .A1(_10309_ ), .A2(_04096_ ), .A3(_04149_ ), .A4(_04155_ ), .ZN(_04180_ ) );
OAI21_X1 _18497_ ( .A(\u_lsu.pmem[2819] ), .B1(_04080_ ), .B2(_11224_ ), .ZN(_04181_ ) );
AOI21_X1 _18498_ ( .A(fanout_net_52 ), .B1(_04180_ ), .B2(_04181_ ), .ZN(_01514_ ) );
BUF_X4 _18499_ ( .A(_03396_ ), .Z(_04182_ ) );
NAND4_X1 _18500_ ( .A1(_03970_ ), .A2(_04182_ ), .A3(_04149_ ), .A4(_10313_ ), .ZN(_04183_ ) );
OAI21_X1 _18501_ ( .A(\u_lsu.pmem[2818] ), .B1(_04080_ ), .B2(_11224_ ), .ZN(_04184_ ) );
AOI21_X1 _18502_ ( .A(fanout_net_52 ), .B1(_04183_ ), .B2(_04184_ ), .ZN(_01515_ ) );
BUF_X4 _18503_ ( .A(_03875_ ), .Z(_04185_ ) );
NAND4_X1 _18504_ ( .A1(_10316_ ), .A2(_04182_ ), .A3(_04185_ ), .A4(_04155_ ), .ZN(_04186_ ) );
BUF_X4 _18505_ ( .A(_03919_ ), .Z(_04187_ ) );
OAI21_X1 _18506_ ( .A(\u_lsu.pmem[2817] ), .B1(_04187_ ), .B2(_11224_ ), .ZN(_04188_ ) );
AOI21_X1 _18507_ ( .A(fanout_net_52 ), .B1(_04186_ ), .B2(_04188_ ), .ZN(_01516_ ) );
NAND4_X1 _18508_ ( .A1(_10320_ ), .A2(_04182_ ), .A3(_04185_ ), .A4(_04155_ ), .ZN(_04189_ ) );
OAI21_X1 _18509_ ( .A(\u_lsu.pmem[2816] ), .B1(_04187_ ), .B2(_11224_ ), .ZN(_04190_ ) );
AOI21_X1 _18510_ ( .A(fanout_net_53 ), .B1(_04189_ ), .B2(_04190_ ), .ZN(_01517_ ) );
NOR2_X1 _18511_ ( .A1(_03850_ ), .A2(_11246_ ), .ZN(_04191_ ) );
NOR2_X1 _18512_ ( .A1(_04191_ ), .A2(\u_lsu.pmem[2791] ), .ZN(_04192_ ) );
AOI211_X1 _18513_ ( .A(fanout_net_53 ), .B(_04192_ ), .C1(_09568_ ), .C2(_04191_ ), .ZN(_01518_ ) );
NAND4_X1 _18514_ ( .A1(_10332_ ), .A2(_04182_ ), .A3(_04185_ ), .A4(_04155_ ), .ZN(_04193_ ) );
OAI21_X1 _18515_ ( .A(\u_lsu.pmem[2790] ), .B1(_04187_ ), .B2(_11247_ ), .ZN(_04194_ ) );
AOI21_X1 _18516_ ( .A(fanout_net_53 ), .B1(_04193_ ), .B2(_04194_ ), .ZN(_01519_ ) );
BUF_X4 _18517_ ( .A(_04154_ ), .Z(_04195_ ) );
NAND4_X1 _18518_ ( .A1(_10336_ ), .A2(_04182_ ), .A3(_04185_ ), .A4(_04195_ ), .ZN(_04196_ ) );
OAI21_X1 _18519_ ( .A(\u_lsu.pmem[2789] ), .B1(_04187_ ), .B2(_11247_ ), .ZN(_04197_ ) );
AOI21_X1 _18520_ ( .A(fanout_net_53 ), .B1(_04196_ ), .B2(_04197_ ), .ZN(_01520_ ) );
NAND4_X1 _18521_ ( .A1(_09703_ ), .A2(_04182_ ), .A3(_03886_ ), .A4(_04097_ ), .ZN(_04198_ ) );
OAI21_X1 _18522_ ( .A(\u_lsu.pmem[4384] ), .B1(_09440_ ), .B2(_09516_ ), .ZN(_04199_ ) );
AOI21_X1 _18523_ ( .A(fanout_net_53 ), .B1(_04198_ ), .B2(_04199_ ), .ZN(_01521_ ) );
OAI21_X1 _18524_ ( .A(\u_lsu.pmem[4228] ), .B1(_09890_ ), .B2(_09882_ ), .ZN(_04200_ ) );
NAND4_X1 _18525_ ( .A1(_02301_ ), .A2(_03064_ ), .A3(_03640_ ), .A4(_03646_ ), .ZN(_04201_ ) );
AOI21_X1 _18526_ ( .A(fanout_net_53 ), .B1(_04200_ ), .B2(_04201_ ), .ZN(_01522_ ) );
NAND4_X1 _18527_ ( .A1(_10339_ ), .A2(_04182_ ), .A3(_04185_ ), .A4(_04195_ ), .ZN(_04202_ ) );
OAI21_X1 _18528_ ( .A(\u_lsu.pmem[2788] ), .B1(_04187_ ), .B2(_11246_ ), .ZN(_04203_ ) );
AOI21_X1 _18529_ ( .A(fanout_net_53 ), .B1(_04202_ ), .B2(_04203_ ), .ZN(_01523_ ) );
NAND4_X1 _18530_ ( .A1(_10345_ ), .A2(_04182_ ), .A3(_04185_ ), .A4(_04195_ ), .ZN(_04204_ ) );
OAI21_X1 _18531_ ( .A(\u_lsu.pmem[2787] ), .B1(_04187_ ), .B2(_11246_ ), .ZN(_04205_ ) );
AOI21_X1 _18532_ ( .A(fanout_net_53 ), .B1(_04204_ ), .B2(_04205_ ), .ZN(_01524_ ) );
NAND4_X1 _18533_ ( .A1(_10350_ ), .A2(_04182_ ), .A3(_04185_ ), .A4(_04195_ ), .ZN(_04206_ ) );
OAI21_X1 _18534_ ( .A(\u_lsu.pmem[2786] ), .B1(_04187_ ), .B2(_11246_ ), .ZN(_04207_ ) );
AOI21_X1 _18535_ ( .A(fanout_net_53 ), .B1(_04206_ ), .B2(_04207_ ), .ZN(_01525_ ) );
NAND4_X1 _18536_ ( .A1(_10354_ ), .A2(_04182_ ), .A3(_04185_ ), .A4(_04195_ ), .ZN(_04208_ ) );
OAI21_X1 _18537_ ( .A(\u_lsu.pmem[2785] ), .B1(_04187_ ), .B2(_11246_ ), .ZN(_04209_ ) );
AOI21_X1 _18538_ ( .A(fanout_net_53 ), .B1(_04208_ ), .B2(_04209_ ), .ZN(_01526_ ) );
BUF_X8 _18539_ ( .A(_09539_ ), .Z(_04210_ ) );
BUF_X4 _18540_ ( .A(_04210_ ), .Z(_04211_ ) );
NAND4_X1 _18541_ ( .A1(_10357_ ), .A2(_04211_ ), .A3(_04185_ ), .A4(_04195_ ), .ZN(_04212_ ) );
OAI21_X1 _18542_ ( .A(\u_lsu.pmem[2784] ), .B1(_04187_ ), .B2(_11246_ ), .ZN(_04213_ ) );
AOI21_X1 _18543_ ( .A(fanout_net_53 ), .B1(_04212_ ), .B2(_04213_ ), .ZN(_01527_ ) );
NOR2_X1 _18544_ ( .A1(_03850_ ), .A2(_11268_ ), .ZN(_04214_ ) );
NOR2_X1 _18545_ ( .A1(_04214_ ), .A2(\u_lsu.pmem[2759] ), .ZN(_04215_ ) );
BUF_X4 _18546_ ( .A(_09567_ ), .Z(_04216_ ) );
AOI211_X1 _18547_ ( .A(fanout_net_53 ), .B(_04215_ ), .C1(_04216_ ), .C2(_04214_ ), .ZN(_01528_ ) );
NAND4_X1 _18548_ ( .A1(_10368_ ), .A2(_04211_ ), .A3(_04185_ ), .A4(_04195_ ), .ZN(_04217_ ) );
OAI21_X1 _18549_ ( .A(\u_lsu.pmem[2758] ), .B1(_04187_ ), .B2(_11269_ ), .ZN(_04218_ ) );
AOI21_X1 _18550_ ( .A(fanout_net_53 ), .B1(_04217_ ), .B2(_04218_ ), .ZN(_01529_ ) );
BUF_X4 _18551_ ( .A(_03875_ ), .Z(_04219_ ) );
NAND4_X1 _18552_ ( .A1(_10371_ ), .A2(_04211_ ), .A3(_04219_ ), .A4(_04195_ ), .ZN(_04220_ ) );
BUF_X4 _18553_ ( .A(_03919_ ), .Z(_04221_ ) );
OAI21_X1 _18554_ ( .A(\u_lsu.pmem[2757] ), .B1(_04221_ ), .B2(_11269_ ), .ZN(_04222_ ) );
AOI21_X1 _18555_ ( .A(fanout_net_53 ), .B1(_04220_ ), .B2(_04222_ ), .ZN(_01530_ ) );
NAND4_X1 _18556_ ( .A1(_10374_ ), .A2(_04211_ ), .A3(_04219_ ), .A4(_04195_ ), .ZN(_04223_ ) );
OAI21_X1 _18557_ ( .A(\u_lsu.pmem[2756] ), .B1(_04221_ ), .B2(_11268_ ), .ZN(_04224_ ) );
AOI21_X1 _18558_ ( .A(fanout_net_53 ), .B1(_04223_ ), .B2(_04224_ ), .ZN(_01531_ ) );
NAND4_X1 _18559_ ( .A1(_10377_ ), .A2(_04211_ ), .A3(_04219_ ), .A4(_04195_ ), .ZN(_04225_ ) );
OAI21_X1 _18560_ ( .A(\u_lsu.pmem[2755] ), .B1(_04221_ ), .B2(_11268_ ), .ZN(_04226_ ) );
AOI21_X1 _18561_ ( .A(fanout_net_53 ), .B1(_04225_ ), .B2(_04226_ ), .ZN(_01532_ ) );
OAI21_X1 _18562_ ( .A(\u_lsu.pmem[4227] ), .B1(_09890_ ), .B2(_09882_ ), .ZN(_04227_ ) );
NAND4_X1 _18563_ ( .A1(_02301_ ), .A2(_09519_ ), .A3(_03640_ ), .A4(_03646_ ), .ZN(_04228_ ) );
AOI21_X1 _18564_ ( .A(fanout_net_53 ), .B1(_04227_ ), .B2(_04228_ ), .ZN(_01533_ ) );
BUF_X4 _18565_ ( .A(_04154_ ), .Z(_04229_ ) );
NAND4_X1 _18566_ ( .A1(_10381_ ), .A2(_04211_ ), .A3(_04219_ ), .A4(_04229_ ), .ZN(_04230_ ) );
OAI21_X1 _18567_ ( .A(\u_lsu.pmem[2754] ), .B1(_04221_ ), .B2(_11268_ ), .ZN(_04231_ ) );
AOI21_X1 _18568_ ( .A(fanout_net_53 ), .B1(_04230_ ), .B2(_04231_ ), .ZN(_01534_ ) );
NAND4_X1 _18569_ ( .A1(_10384_ ), .A2(_04211_ ), .A3(_04219_ ), .A4(_04229_ ), .ZN(_04232_ ) );
OAI21_X1 _18570_ ( .A(\u_lsu.pmem[2753] ), .B1(_04221_ ), .B2(_11268_ ), .ZN(_04233_ ) );
AOI21_X1 _18571_ ( .A(fanout_net_53 ), .B1(_04232_ ), .B2(_04233_ ), .ZN(_01535_ ) );
NAND4_X1 _18572_ ( .A1(_10391_ ), .A2(_04211_ ), .A3(_04219_ ), .A4(_04229_ ), .ZN(_04234_ ) );
OAI21_X1 _18573_ ( .A(\u_lsu.pmem[2752] ), .B1(_04221_ ), .B2(_11268_ ), .ZN(_04235_ ) );
AOI21_X1 _18574_ ( .A(fanout_net_53 ), .B1(_04234_ ), .B2(_04235_ ), .ZN(_01536_ ) );
NAND4_X1 _18575_ ( .A1(_10394_ ), .A2(_04211_ ), .A3(_04219_ ), .A4(_04229_ ), .ZN(_04236_ ) );
BUF_X4 _18576_ ( .A(_09730_ ), .Z(_04237_ ) );
OAI21_X1 _18577_ ( .A(\u_lsu.pmem[2727] ), .B1(_11294_ ), .B2(_04237_ ), .ZN(_04238_ ) );
AOI21_X1 _18578_ ( .A(fanout_net_53 ), .B1(_04236_ ), .B2(_04238_ ), .ZN(_01537_ ) );
NAND4_X1 _18579_ ( .A1(_10402_ ), .A2(_04211_ ), .A3(_04219_ ), .A4(_04229_ ), .ZN(_04239_ ) );
OAI21_X1 _18580_ ( .A(\u_lsu.pmem[2726] ), .B1(_11294_ ), .B2(_04237_ ), .ZN(_04240_ ) );
AOI21_X1 _18581_ ( .A(fanout_net_53 ), .B1(_04239_ ), .B2(_04240_ ), .ZN(_01538_ ) );
BUF_X4 _18582_ ( .A(_04210_ ), .Z(_04241_ ) );
NAND4_X1 _18583_ ( .A1(_10405_ ), .A2(_04241_ ), .A3(_04219_ ), .A4(_04229_ ), .ZN(_04242_ ) );
OAI21_X1 _18584_ ( .A(\u_lsu.pmem[2725] ), .B1(_11294_ ), .B2(_04237_ ), .ZN(_04243_ ) );
AOI21_X1 _18585_ ( .A(fanout_net_53 ), .B1(_04242_ ), .B2(_04243_ ), .ZN(_01539_ ) );
NAND4_X1 _18586_ ( .A1(_10408_ ), .A2(_04241_ ), .A3(_04219_ ), .A4(_04229_ ), .ZN(_04244_ ) );
OAI21_X1 _18587_ ( .A(\u_lsu.pmem[2724] ), .B1(_11294_ ), .B2(_04237_ ), .ZN(_04245_ ) );
AOI21_X1 _18588_ ( .A(fanout_net_53 ), .B1(_04244_ ), .B2(_04245_ ), .ZN(_01540_ ) );
BUF_X4 _18589_ ( .A(_03875_ ), .Z(_04246_ ) );
NAND4_X1 _18590_ ( .A1(_10411_ ), .A2(_04241_ ), .A3(_04246_ ), .A4(_04229_ ), .ZN(_04247_ ) );
OAI21_X1 _18591_ ( .A(\u_lsu.pmem[2723] ), .B1(_11294_ ), .B2(_04237_ ), .ZN(_04248_ ) );
AOI21_X1 _18592_ ( .A(fanout_net_53 ), .B1(_04247_ ), .B2(_04248_ ), .ZN(_01541_ ) );
NAND4_X1 _18593_ ( .A1(_10414_ ), .A2(_04241_ ), .A3(_04246_ ), .A4(_04229_ ), .ZN(_04249_ ) );
OAI21_X1 _18594_ ( .A(\u_lsu.pmem[2722] ), .B1(_11294_ ), .B2(_04237_ ), .ZN(_04250_ ) );
AOI21_X1 _18595_ ( .A(fanout_net_53 ), .B1(_04249_ ), .B2(_04250_ ), .ZN(_01542_ ) );
NAND4_X1 _18596_ ( .A1(_10417_ ), .A2(_04241_ ), .A3(_04246_ ), .A4(_04229_ ), .ZN(_04251_ ) );
OAI21_X1 _18597_ ( .A(\u_lsu.pmem[2721] ), .B1(_11294_ ), .B2(_04237_ ), .ZN(_04252_ ) );
AOI21_X1 _18598_ ( .A(fanout_net_53 ), .B1(_04251_ ), .B2(_04252_ ), .ZN(_01543_ ) );
OAI21_X1 _18599_ ( .A(\u_lsu.pmem[4226] ), .B1(_09890_ ), .B2(_09882_ ), .ZN(_04253_ ) );
NAND4_X1 _18600_ ( .A1(_09906_ ), .A2(_03361_ ), .A3(_03640_ ), .A4(_03646_ ), .ZN(_04254_ ) );
AOI21_X1 _18601_ ( .A(fanout_net_53 ), .B1(_04253_ ), .B2(_04254_ ), .ZN(_01544_ ) );
NAND4_X1 _18602_ ( .A1(_03970_ ), .A2(_02935_ ), .A3(_03753_ ), .A4(_11292_ ), .ZN(_04255_ ) );
OAI21_X1 _18603_ ( .A(\u_lsu.pmem[2720] ), .B1(_11294_ ), .B2(_04237_ ), .ZN(_04256_ ) );
AOI21_X1 _18604_ ( .A(fanout_net_53 ), .B1(_04255_ ), .B2(_04256_ ), .ZN(_01545_ ) );
OAI21_X1 _18605_ ( .A(\u_lsu.pmem[2695] ), .B1(_11317_ ), .B2(_04163_ ), .ZN(_04257_ ) );
NAND4_X1 _18606_ ( .A1(_10436_ ), .A2(_03361_ ), .A3(_04093_ ), .A4(_04094_ ), .ZN(_04258_ ) );
AOI21_X1 _18607_ ( .A(fanout_net_53 ), .B1(_04257_ ), .B2(_04258_ ), .ZN(_01546_ ) );
BUF_X4 _18608_ ( .A(_04154_ ), .Z(_04259_ ) );
NAND4_X1 _18609_ ( .A1(_03457_ ), .A2(_09658_ ), .A3(_04246_ ), .A4(_04259_ ), .ZN(_04260_ ) );
OAI21_X1 _18610_ ( .A(\u_lsu.pmem[2694] ), .B1(_11316_ ), .B2(_04237_ ), .ZN(_04261_ ) );
AOI21_X1 _18611_ ( .A(fanout_net_54 ), .B1(_04260_ ), .B2(_04261_ ), .ZN(_01547_ ) );
NAND4_X1 _18612_ ( .A1(_03457_ ), .A2(_09713_ ), .A3(_04246_ ), .A4(_04259_ ), .ZN(_04262_ ) );
OAI21_X1 _18613_ ( .A(\u_lsu.pmem[2693] ), .B1(_11316_ ), .B2(_04237_ ), .ZN(_04263_ ) );
AOI21_X1 _18614_ ( .A(fanout_net_54 ), .B1(_04262_ ), .B2(_04263_ ), .ZN(_01548_ ) );
NAND4_X1 _18615_ ( .A1(_03457_ ), .A2(_09514_ ), .A3(_04246_ ), .A4(_04259_ ), .ZN(_04264_ ) );
BUF_X8 _18616_ ( .A(_09450_ ), .Z(_04265_ ) );
BUF_X4 _18617_ ( .A(_04265_ ), .Z(_04266_ ) );
OAI21_X1 _18618_ ( .A(\u_lsu.pmem[2692] ), .B1(_11316_ ), .B2(_04266_ ), .ZN(_04267_ ) );
AOI21_X1 _18619_ ( .A(fanout_net_54 ), .B1(_04264_ ), .B2(_04267_ ), .ZN(_01549_ ) );
NAND4_X1 _18620_ ( .A1(_03457_ ), .A2(_10456_ ), .A3(_04246_ ), .A4(_04259_ ), .ZN(_04268_ ) );
OAI21_X1 _18621_ ( .A(\u_lsu.pmem[2691] ), .B1(_11316_ ), .B2(_04266_ ), .ZN(_04269_ ) );
AOI21_X1 _18622_ ( .A(fanout_net_54 ), .B1(_04268_ ), .B2(_04269_ ), .ZN(_01550_ ) );
OAI21_X1 _18623_ ( .A(\u_lsu.pmem[2690] ), .B1(_11317_ ), .B2(_04163_ ), .ZN(_04270_ ) );
NAND4_X1 _18624_ ( .A1(_10460_ ), .A2(_03361_ ), .A3(_04093_ ), .A4(_04094_ ), .ZN(_04271_ ) );
AOI21_X1 _18625_ ( .A(fanout_net_54 ), .B1(_04270_ ), .B2(_04271_ ), .ZN(_01551_ ) );
NAND4_X1 _18626_ ( .A1(_03457_ ), .A2(_09544_ ), .A3(_04246_ ), .A4(_04259_ ), .ZN(_04272_ ) );
OAI21_X1 _18627_ ( .A(\u_lsu.pmem[2689] ), .B1(_11316_ ), .B2(_04266_ ), .ZN(_04273_ ) );
AOI21_X1 _18628_ ( .A(fanout_net_54 ), .B1(_04272_ ), .B2(_04273_ ), .ZN(_01552_ ) );
NAND4_X1 _18629_ ( .A1(_03457_ ), .A2(_10467_ ), .A3(_04246_ ), .A4(_04259_ ), .ZN(_04274_ ) );
OAI21_X1 _18630_ ( .A(\u_lsu.pmem[2688] ), .B1(_11316_ ), .B2(_04266_ ), .ZN(_04275_ ) );
AOI21_X1 _18631_ ( .A(fanout_net_54 ), .B1(_04274_ ), .B2(_04275_ ), .ZN(_01553_ ) );
NOR2_X4 _18632_ ( .A1(_09450_ ), .A2(_11342_ ), .ZN(_04276_ ) );
NOR2_X1 _18633_ ( .A1(_04276_ ), .A2(\u_lsu.pmem[2663] ), .ZN(_04277_ ) );
AOI211_X1 _18634_ ( .A(fanout_net_54 ), .B(_04277_ ), .C1(_04216_ ), .C2(_04276_ ), .ZN(_01554_ ) );
OAI21_X1 _18635_ ( .A(\u_lsu.pmem[4225] ), .B1(_09890_ ), .B2(_09882_ ), .ZN(_04278_ ) );
BUF_X4 _18636_ ( .A(_02881_ ), .Z(_04279_ ) );
NAND4_X1 _18637_ ( .A1(_02301_ ), .A2(_02308_ ), .A3(_04279_ ), .A4(_03646_ ), .ZN(_04280_ ) );
AOI21_X1 _18638_ ( .A(fanout_net_54 ), .B1(_04278_ ), .B2(_04280_ ), .ZN(_01555_ ) );
NAND2_X1 _18639_ ( .A1(_04276_ ), .A2(_11145_ ), .ZN(_04281_ ) );
OAI21_X1 _18640_ ( .A(\u_lsu.pmem[2662] ), .B1(_04221_ ), .B2(_11343_ ), .ZN(_04282_ ) );
AOI21_X1 _18641_ ( .A(fanout_net_54 ), .B1(_04281_ ), .B2(_04282_ ), .ZN(_01556_ ) );
NAND2_X1 _18642_ ( .A1(_04276_ ), .A2(_11148_ ), .ZN(_04283_ ) );
OAI21_X1 _18643_ ( .A(\u_lsu.pmem[2661] ), .B1(_04221_ ), .B2(_11343_ ), .ZN(_04284_ ) );
AOI21_X1 _18644_ ( .A(fanout_net_54 ), .B1(_04283_ ), .B2(_04284_ ), .ZN(_01557_ ) );
NAND2_X1 _18645_ ( .A1(_04276_ ), .A2(_03084_ ), .ZN(_04285_ ) );
OAI21_X1 _18646_ ( .A(\u_lsu.pmem[2660] ), .B1(_04221_ ), .B2(_11342_ ), .ZN(_04286_ ) );
AOI21_X1 _18647_ ( .A(fanout_net_54 ), .B1(_04285_ ), .B2(_04286_ ), .ZN(_01558_ ) );
NAND2_X1 _18648_ ( .A1(_04276_ ), .A2(_03114_ ), .ZN(_04287_ ) );
OAI21_X1 _18649_ ( .A(\u_lsu.pmem[2659] ), .B1(_04221_ ), .B2(_11342_ ), .ZN(_04288_ ) );
AOI21_X1 _18650_ ( .A(fanout_net_54 ), .B1(_04287_ ), .B2(_04288_ ), .ZN(_01559_ ) );
NAND2_X1 _18651_ ( .A1(_04276_ ), .A2(_03145_ ), .ZN(_04289_ ) );
BUF_X4 _18652_ ( .A(_03919_ ), .Z(_04290_ ) );
OAI21_X1 _18653_ ( .A(\u_lsu.pmem[2658] ), .B1(_04290_ ), .B2(_11342_ ), .ZN(_04291_ ) );
AOI21_X1 _18654_ ( .A(fanout_net_54 ), .B1(_04289_ ), .B2(_04291_ ), .ZN(_01560_ ) );
NAND2_X1 _18655_ ( .A1(_04276_ ), .A2(_03174_ ), .ZN(_04292_ ) );
OAI21_X1 _18656_ ( .A(\u_lsu.pmem[2657] ), .B1(_04290_ ), .B2(_11342_ ), .ZN(_04293_ ) );
AOI21_X1 _18657_ ( .A(fanout_net_54 ), .B1(_04292_ ), .B2(_04293_ ), .ZN(_01561_ ) );
NAND2_X1 _18658_ ( .A1(_04276_ ), .A2(_03203_ ), .ZN(_04294_ ) );
OAI21_X1 _18659_ ( .A(\u_lsu.pmem[2656] ), .B1(_04290_ ), .B2(_11342_ ), .ZN(_04295_ ) );
AOI21_X1 _18660_ ( .A(fanout_net_54 ), .B1(_04294_ ), .B2(_04295_ ), .ZN(_01562_ ) );
BUF_X4 _18661_ ( .A(_09953_ ), .Z(_04296_ ) );
NAND4_X1 _18662_ ( .A1(_04296_ ), .A2(_02935_ ), .A3(_09914_ ), .A4(_11373_ ), .ZN(_04297_ ) );
OAI21_X1 _18663_ ( .A(\u_lsu.pmem[2631] ), .B1(_11371_ ), .B2(_04266_ ), .ZN(_04298_ ) );
AOI21_X1 _18664_ ( .A(fanout_net_54 ), .B1(_04297_ ), .B2(_04298_ ), .ZN(_01563_ ) );
NAND4_X1 _18665_ ( .A1(_04296_ ), .A2(_02935_ ), .A3(_09925_ ), .A4(_11373_ ), .ZN(_04299_ ) );
OAI21_X1 _18666_ ( .A(\u_lsu.pmem[2630] ), .B1(_11371_ ), .B2(_04266_ ), .ZN(_04300_ ) );
AOI21_X1 _18667_ ( .A(fanout_net_54 ), .B1(_04299_ ), .B2(_04300_ ), .ZN(_01564_ ) );
NAND4_X1 _18668_ ( .A1(_04296_ ), .A2(_02935_ ), .A3(_09928_ ), .A4(_11373_ ), .ZN(_04301_ ) );
OAI21_X1 _18669_ ( .A(\u_lsu.pmem[2629] ), .B1(_11371_ ), .B2(_04266_ ), .ZN(_04302_ ) );
AOI21_X1 _18670_ ( .A(fanout_net_54 ), .B1(_04301_ ), .B2(_04302_ ), .ZN(_01565_ ) );
OAI21_X1 _18671_ ( .A(\u_lsu.pmem[4224] ), .B1(_09890_ ), .B2(_09882_ ), .ZN(_04303_ ) );
NAND4_X1 _18672_ ( .A1(_09893_ ), .A2(_09547_ ), .A3(_04279_ ), .A4(_03646_ ), .ZN(_04304_ ) );
AOI21_X1 _18673_ ( .A(fanout_net_54 ), .B1(_04303_ ), .B2(_04304_ ), .ZN(_01566_ ) );
NAND4_X1 _18674_ ( .A1(_04296_ ), .A2(_10066_ ), .A3(_11151_ ), .A4(_11373_ ), .ZN(_04305_ ) );
OAI21_X1 _18675_ ( .A(\u_lsu.pmem[2628] ), .B1(_11371_ ), .B2(_04266_ ), .ZN(_04306_ ) );
AOI21_X1 _18676_ ( .A(fanout_net_54 ), .B1(_04305_ ), .B2(_04306_ ), .ZN(_01567_ ) );
NAND4_X1 _18677_ ( .A1(_04296_ ), .A2(_10066_ ), .A3(_09934_ ), .A4(_11373_ ), .ZN(_04307_ ) );
OAI21_X1 _18678_ ( .A(\u_lsu.pmem[2627] ), .B1(_11371_ ), .B2(_04266_ ), .ZN(_04308_ ) );
AOI21_X1 _18679_ ( .A(fanout_net_54 ), .B1(_04307_ ), .B2(_04308_ ), .ZN(_01568_ ) );
NAND4_X1 _18680_ ( .A1(_04296_ ), .A2(_10066_ ), .A3(_10015_ ), .A4(_11373_ ), .ZN(_04309_ ) );
OAI21_X1 _18681_ ( .A(\u_lsu.pmem[2626] ), .B1(_11371_ ), .B2(_04266_ ), .ZN(_04310_ ) );
AOI21_X1 _18682_ ( .A(fanout_net_54 ), .B1(_04309_ ), .B2(_04310_ ), .ZN(_01569_ ) );
NAND4_X1 _18683_ ( .A1(_04296_ ), .A2(_10066_ ), .A3(_09941_ ), .A4(_11373_ ), .ZN(_04311_ ) );
BUF_X4 _18684_ ( .A(_04265_ ), .Z(_04312_ ) );
OAI21_X1 _18685_ ( .A(\u_lsu.pmem[2625] ), .B1(_11371_ ), .B2(_04312_ ), .ZN(_04313_ ) );
AOI21_X1 _18686_ ( .A(fanout_net_54 ), .B1(_04311_ ), .B2(_04313_ ), .ZN(_01570_ ) );
NAND4_X1 _18687_ ( .A1(_04296_ ), .A2(_10066_ ), .A3(_03753_ ), .A4(_11373_ ), .ZN(_04314_ ) );
OAI21_X1 _18688_ ( .A(\u_lsu.pmem[2624] ), .B1(_11371_ ), .B2(_04312_ ), .ZN(_04315_ ) );
AOI21_X1 _18689_ ( .A(fanout_net_54 ), .B1(_04314_ ), .B2(_04315_ ), .ZN(_01571_ ) );
NAND4_X1 _18690_ ( .A1(_10527_ ), .A2(_04241_ ), .A3(_04246_ ), .A4(_04259_ ), .ZN(_04316_ ) );
OAI21_X1 _18691_ ( .A(\u_lsu.pmem[2599] ), .B1(_04290_ ), .B2(_11398_ ), .ZN(_04317_ ) );
AOI21_X1 _18692_ ( .A(fanout_net_54 ), .B1(_04316_ ), .B2(_04317_ ), .ZN(_01572_ ) );
BUF_X4 _18693_ ( .A(_03875_ ), .Z(_04318_ ) );
NAND4_X1 _18694_ ( .A1(_10535_ ), .A2(_04241_ ), .A3(_04318_ ), .A4(_04259_ ), .ZN(_04319_ ) );
OAI21_X1 _18695_ ( .A(\u_lsu.pmem[2598] ), .B1(_04290_ ), .B2(_11398_ ), .ZN(_04320_ ) );
AOI21_X1 _18696_ ( .A(fanout_net_54 ), .B1(_04319_ ), .B2(_04320_ ), .ZN(_01573_ ) );
NAND4_X1 _18697_ ( .A1(_10538_ ), .A2(_04241_ ), .A3(_04318_ ), .A4(_04259_ ), .ZN(_04321_ ) );
OAI21_X1 _18698_ ( .A(\u_lsu.pmem[2597] ), .B1(_04290_ ), .B2(_11397_ ), .ZN(_04322_ ) );
AOI21_X1 _18699_ ( .A(fanout_net_54 ), .B1(_04321_ ), .B2(_04322_ ), .ZN(_01574_ ) );
NOR2_X2 _18700_ ( .A1(_09141_ ), .A2(_11397_ ), .ZN(_04323_ ) );
OAI21_X1 _18701_ ( .A(_09109_ ), .B1(_04323_ ), .B2(\u_lsu.pmem[2596] ), .ZN(_04324_ ) );
AOI21_X1 _18702_ ( .A(_04324_ ), .B1(_09691_ ), .B2(_04323_ ), .ZN(_01575_ ) );
NAND2_X1 _18703_ ( .A1(_04323_ ), .A2(_03114_ ), .ZN(_04325_ ) );
OAI21_X1 _18704_ ( .A(\u_lsu.pmem[2595] ), .B1(_04290_ ), .B2(_11397_ ), .ZN(_04326_ ) );
AOI21_X1 _18705_ ( .A(fanout_net_54 ), .B1(_04325_ ), .B2(_04326_ ), .ZN(_01576_ ) );
OAI21_X1 _18706_ ( .A(\u_lsu.pmem[4199] ), .B1(_03705_ ), .B2(_09920_ ), .ZN(_04327_ ) );
NAND4_X1 _18707_ ( .A1(_09742_ ), .A2(_03504_ ), .A3(_04279_ ), .A4(_02323_ ), .ZN(_04328_ ) );
AOI21_X1 _18708_ ( .A(fanout_net_54 ), .B1(_04327_ ), .B2(_04328_ ), .ZN(_01577_ ) );
NAND2_X1 _18709_ ( .A1(_04323_ ), .A2(_03145_ ), .ZN(_04329_ ) );
OAI21_X1 _18710_ ( .A(\u_lsu.pmem[2594] ), .B1(_04290_ ), .B2(_11397_ ), .ZN(_04330_ ) );
AOI21_X1 _18711_ ( .A(fanout_net_55 ), .B1(_04329_ ), .B2(_04330_ ), .ZN(_01578_ ) );
NAND2_X1 _18712_ ( .A1(_04323_ ), .A2(_03174_ ), .ZN(_04331_ ) );
OAI21_X1 _18713_ ( .A(\u_lsu.pmem[2593] ), .B1(_04290_ ), .B2(_11397_ ), .ZN(_04332_ ) );
AOI21_X1 _18714_ ( .A(fanout_net_55 ), .B1(_04331_ ), .B2(_04332_ ), .ZN(_01579_ ) );
NAND4_X1 _18715_ ( .A1(_10556_ ), .A2(_04241_ ), .A3(_04318_ ), .A4(_04259_ ), .ZN(_04333_ ) );
OAI21_X1 _18716_ ( .A(\u_lsu.pmem[2592] ), .B1(_04290_ ), .B2(_11397_ ), .ZN(_04334_ ) );
AOI21_X1 _18717_ ( .A(fanout_net_55 ), .B1(_04333_ ), .B2(_04334_ ), .ZN(_01580_ ) );
OAI21_X1 _18718_ ( .A(\u_lsu.pmem[2567] ), .B1(_11420_ ), .B2(_04163_ ), .ZN(_04335_ ) );
NAND3_X1 _18719_ ( .A1(_04161_ ), .A2(_11423_ ), .A3(_11422_ ), .ZN(_04336_ ) );
AOI21_X1 _18720_ ( .A(fanout_net_55 ), .B1(_04335_ ), .B2(_04336_ ), .ZN(_01581_ ) );
OAI21_X1 _18721_ ( .A(\u_lsu.pmem[2566] ), .B1(_11420_ ), .B2(_04163_ ), .ZN(_04337_ ) );
NAND3_X1 _18722_ ( .A1(_04161_ ), .A2(_10444_ ), .A3(_11422_ ), .ZN(_04338_ ) );
AOI21_X1 _18723_ ( .A(fanout_net_55 ), .B1(_04337_ ), .B2(_04338_ ), .ZN(_01582_ ) );
OAI21_X1 _18724_ ( .A(\u_lsu.pmem[2565] ), .B1(_11420_ ), .B2(_04163_ ), .ZN(_04339_ ) );
NAND3_X1 _18725_ ( .A1(_04161_ ), .A2(_10448_ ), .A3(_11422_ ), .ZN(_04340_ ) );
AOI21_X1 _18726_ ( .A(fanout_net_55 ), .B1(_04339_ ), .B2(_04340_ ), .ZN(_01583_ ) );
OAI21_X1 _18727_ ( .A(\u_lsu.pmem[2564] ), .B1(_11420_ ), .B2(_04163_ ), .ZN(_04341_ ) );
NAND3_X1 _18728_ ( .A1(_04161_ ), .A2(_10453_ ), .A3(_11422_ ), .ZN(_04342_ ) );
AOI21_X1 _18729_ ( .A(fanout_net_55 ), .B1(_04341_ ), .B2(_04342_ ), .ZN(_01584_ ) );
NAND4_X1 _18730_ ( .A1(_10575_ ), .A2(_09882_ ), .A3(_09979_ ), .A4(_03978_ ), .ZN(_04343_ ) );
OAI21_X1 _18731_ ( .A(\u_lsu.pmem[2563] ), .B1(_11419_ ), .B2(_04312_ ), .ZN(_04344_ ) );
AOI21_X1 _18732_ ( .A(fanout_net_55 ), .B1(_04343_ ), .B2(_04344_ ), .ZN(_01585_ ) );
BUF_X4 _18733_ ( .A(_04154_ ), .Z(_04345_ ) );
NAND4_X1 _18734_ ( .A1(_10584_ ), .A2(_09806_ ), .A3(_04318_ ), .A4(_04345_ ), .ZN(_04346_ ) );
OAI21_X1 _18735_ ( .A(\u_lsu.pmem[2562] ), .B1(_11419_ ), .B2(_04312_ ), .ZN(_04347_ ) );
AOI21_X1 _18736_ ( .A(fanout_net_55 ), .B1(_04346_ ), .B2(_04347_ ), .ZN(_01586_ ) );
OAI21_X1 _18737_ ( .A(\u_lsu.pmem[2561] ), .B1(_11420_ ), .B2(_04163_ ), .ZN(_04348_ ) );
NAND3_X1 _18738_ ( .A1(_04161_ ), .A2(_10463_ ), .A3(_11422_ ), .ZN(_04349_ ) );
AOI21_X1 _18739_ ( .A(fanout_net_55 ), .B1(_04348_ ), .B2(_04349_ ), .ZN(_01587_ ) );
OAI21_X1 _18740_ ( .A(\u_lsu.pmem[4198] ), .B1(_03705_ ), .B2(_09920_ ), .ZN(_04350_ ) );
NAND4_X1 _18741_ ( .A1(_11347_ ), .A2(_03504_ ), .A3(_04279_ ), .A4(_02323_ ), .ZN(_04351_ ) );
AOI21_X1 _18742_ ( .A(fanout_net_55 ), .B1(_04350_ ), .B2(_04351_ ), .ZN(_01588_ ) );
NAND4_X1 _18743_ ( .A1(_10591_ ), .A2(_09676_ ), .A3(_09979_ ), .A4(_03978_ ), .ZN(_04352_ ) );
OAI21_X1 _18744_ ( .A(\u_lsu.pmem[2560] ), .B1(_11419_ ), .B2(_04312_ ), .ZN(_04353_ ) );
AOI21_X1 _18745_ ( .A(fanout_net_55 ), .B1(_04352_ ), .B2(_04353_ ), .ZN(_01589_ ) );
NOR2_X2 _18746_ ( .A1(_03850_ ), .A2(_11443_ ), .ZN(_04354_ ) );
NOR2_X1 _18747_ ( .A1(_04354_ ), .A2(\u_lsu.pmem[2535] ), .ZN(_04355_ ) );
AOI211_X1 _18748_ ( .A(fanout_net_55 ), .B(_04355_ ), .C1(_04216_ ), .C2(_04354_ ), .ZN(_01590_ ) );
NAND4_X1 _18749_ ( .A1(_10603_ ), .A2(_04241_ ), .A3(_04318_ ), .A4(_04345_ ), .ZN(_04356_ ) );
BUF_X4 _18750_ ( .A(_03919_ ), .Z(_04357_ ) );
OAI21_X1 _18751_ ( .A(\u_lsu.pmem[2534] ), .B1(_04357_ ), .B2(_11444_ ), .ZN(_04358_ ) );
AOI21_X1 _18752_ ( .A(fanout_net_55 ), .B1(_04356_ ), .B2(_04358_ ), .ZN(_01591_ ) );
BUF_X4 _18753_ ( .A(_04210_ ), .Z(_04359_ ) );
NAND4_X1 _18754_ ( .A1(_10608_ ), .A2(_04359_ ), .A3(_04318_ ), .A4(_04345_ ), .ZN(_04360_ ) );
OAI21_X1 _18755_ ( .A(\u_lsu.pmem[2533] ), .B1(_04357_ ), .B2(_11444_ ), .ZN(_04361_ ) );
AOI21_X1 _18756_ ( .A(fanout_net_55 ), .B1(_04360_ ), .B2(_04361_ ), .ZN(_01592_ ) );
NAND4_X1 _18757_ ( .A1(_10611_ ), .A2(_04359_ ), .A3(_04318_ ), .A4(_04345_ ), .ZN(_04362_ ) );
OAI21_X1 _18758_ ( .A(\u_lsu.pmem[2532] ), .B1(_04357_ ), .B2(_11443_ ), .ZN(_04363_ ) );
AOI21_X1 _18759_ ( .A(fanout_net_55 ), .B1(_04362_ ), .B2(_04363_ ), .ZN(_01593_ ) );
NAND4_X1 _18760_ ( .A1(_10614_ ), .A2(_04359_ ), .A3(_04318_ ), .A4(_04345_ ), .ZN(_04364_ ) );
OAI21_X1 _18761_ ( .A(\u_lsu.pmem[2531] ), .B1(_04357_ ), .B2(_11443_ ), .ZN(_04365_ ) );
AOI21_X1 _18762_ ( .A(fanout_net_55 ), .B1(_04364_ ), .B2(_04365_ ), .ZN(_01594_ ) );
NAND4_X1 _18763_ ( .A1(_10617_ ), .A2(_04359_ ), .A3(_04318_ ), .A4(_04345_ ), .ZN(_04366_ ) );
OAI21_X1 _18764_ ( .A(\u_lsu.pmem[2530] ), .B1(_04357_ ), .B2(_11443_ ), .ZN(_04367_ ) );
AOI21_X1 _18765_ ( .A(fanout_net_55 ), .B1(_04366_ ), .B2(_04367_ ), .ZN(_01595_ ) );
NAND4_X1 _18766_ ( .A1(_10621_ ), .A2(_04359_ ), .A3(_04318_ ), .A4(_04345_ ), .ZN(_04368_ ) );
OAI21_X1 _18767_ ( .A(\u_lsu.pmem[2529] ), .B1(_04357_ ), .B2(_11443_ ), .ZN(_04369_ ) );
AOI21_X1 _18768_ ( .A(fanout_net_55 ), .B1(_04368_ ), .B2(_04369_ ), .ZN(_01596_ ) );
BUF_X4 _18769_ ( .A(_03875_ ), .Z(_04370_ ) );
NAND4_X1 _18770_ ( .A1(_10624_ ), .A2(_04359_ ), .A3(_04370_ ), .A4(_04345_ ), .ZN(_04371_ ) );
OAI21_X1 _18771_ ( .A(\u_lsu.pmem[2528] ), .B1(_04357_ ), .B2(_11443_ ), .ZN(_04372_ ) );
AOI21_X1 _18772_ ( .A(fanout_net_55 ), .B1(_04371_ ), .B2(_04372_ ), .ZN(_01597_ ) );
NOR2_X4 _18773_ ( .A1(_03850_ ), .A2(_11470_ ), .ZN(_04373_ ) );
NOR2_X1 _18774_ ( .A1(_04373_ ), .A2(\u_lsu.pmem[2503] ), .ZN(_04374_ ) );
AOI211_X1 _18775_ ( .A(fanout_net_55 ), .B(_04374_ ), .C1(_04216_ ), .C2(_04373_ ), .ZN(_01598_ ) );
OAI21_X1 _18776_ ( .A(\u_lsu.pmem[4197] ), .B1(_03705_ ), .B2(_09919_ ), .ZN(_04375_ ) );
BUF_X4 _18777_ ( .A(_09950_ ), .Z(_04376_ ) );
NAND4_X1 _18778_ ( .A1(_11351_ ), .A2(_04376_ ), .A3(_04279_ ), .A4(_02323_ ), .ZN(_04377_ ) );
AOI21_X1 _18779_ ( .A(fanout_net_55 ), .B1(_04375_ ), .B2(_04377_ ), .ZN(_01599_ ) );
NAND4_X1 _18780_ ( .A1(_10632_ ), .A2(_04359_ ), .A3(_04370_ ), .A4(_04345_ ), .ZN(_04378_ ) );
OAI21_X1 _18781_ ( .A(\u_lsu.pmem[2502] ), .B1(_04357_ ), .B2(_11471_ ), .ZN(_04379_ ) );
AOI21_X1 _18782_ ( .A(fanout_net_55 ), .B1(_04378_ ), .B2(_04379_ ), .ZN(_01600_ ) );
NAND4_X1 _18783_ ( .A1(_10635_ ), .A2(_04359_ ), .A3(_04370_ ), .A4(_04345_ ), .ZN(_04380_ ) );
OAI21_X1 _18784_ ( .A(\u_lsu.pmem[2501] ), .B1(_04357_ ), .B2(_11471_ ), .ZN(_04381_ ) );
AOI21_X1 _18785_ ( .A(fanout_net_55 ), .B1(_04380_ ), .B2(_04381_ ), .ZN(_01601_ ) );
BUF_X4 _18786_ ( .A(_04154_ ), .Z(_04382_ ) );
NAND4_X1 _18787_ ( .A1(_10641_ ), .A2(_04359_ ), .A3(_04370_ ), .A4(_04382_ ), .ZN(_04383_ ) );
OAI21_X1 _18788_ ( .A(\u_lsu.pmem[2500] ), .B1(_04357_ ), .B2(_11470_ ), .ZN(_04384_ ) );
AOI21_X1 _18789_ ( .A(fanout_net_55 ), .B1(_04383_ ), .B2(_04384_ ), .ZN(_01602_ ) );
NAND4_X1 _18790_ ( .A1(_10645_ ), .A2(_04359_ ), .A3(_04370_ ), .A4(_04382_ ), .ZN(_04385_ ) );
BUF_X4 _18791_ ( .A(_03919_ ), .Z(_04386_ ) );
OAI21_X1 _18792_ ( .A(\u_lsu.pmem[2499] ), .B1(_04386_ ), .B2(_11470_ ), .ZN(_04387_ ) );
AOI21_X1 _18793_ ( .A(fanout_net_55 ), .B1(_04385_ ), .B2(_04387_ ), .ZN(_01603_ ) );
BUF_X4 _18794_ ( .A(_04210_ ), .Z(_04388_ ) );
NAND4_X1 _18795_ ( .A1(_10649_ ), .A2(_04388_ ), .A3(_04370_ ), .A4(_04382_ ), .ZN(_04389_ ) );
OAI21_X1 _18796_ ( .A(\u_lsu.pmem[2498] ), .B1(_04386_ ), .B2(_11470_ ), .ZN(_04390_ ) );
AOI21_X1 _18797_ ( .A(fanout_net_55 ), .B1(_04389_ ), .B2(_04390_ ), .ZN(_01604_ ) );
NAND4_X1 _18798_ ( .A1(_10652_ ), .A2(_04388_ ), .A3(_04370_ ), .A4(_04382_ ), .ZN(_04391_ ) );
OAI21_X1 _18799_ ( .A(\u_lsu.pmem[2497] ), .B1(_04386_ ), .B2(_11470_ ), .ZN(_04392_ ) );
AOI21_X1 _18800_ ( .A(fanout_net_55 ), .B1(_04391_ ), .B2(_04392_ ), .ZN(_01605_ ) );
NAND4_X1 _18801_ ( .A1(_10655_ ), .A2(_04388_ ), .A3(_04370_ ), .A4(_04382_ ), .ZN(_04393_ ) );
OAI21_X1 _18802_ ( .A(\u_lsu.pmem[2496] ), .B1(_04386_ ), .B2(_11470_ ), .ZN(_04394_ ) );
AOI21_X1 _18803_ ( .A(fanout_net_55 ), .B1(_04393_ ), .B2(_04394_ ), .ZN(_01606_ ) );
NAND4_X1 _18804_ ( .A1(_10658_ ), .A2(_04388_ ), .A3(_04370_ ), .A4(_04382_ ), .ZN(_04395_ ) );
OAI21_X1 _18805_ ( .A(\u_lsu.pmem[2471] ), .B1(_11501_ ), .B2(_04312_ ), .ZN(_04396_ ) );
AOI21_X1 _18806_ ( .A(fanout_net_55 ), .B1(_04395_ ), .B2(_04396_ ), .ZN(_01607_ ) );
NAND4_X1 _18807_ ( .A1(_10665_ ), .A2(_04388_ ), .A3(_04370_ ), .A4(_04382_ ), .ZN(_04397_ ) );
OAI21_X1 _18808_ ( .A(\u_lsu.pmem[2470] ), .B1(_11501_ ), .B2(_04312_ ), .ZN(_04398_ ) );
AOI21_X1 _18809_ ( .A(fanout_net_56 ), .B1(_04397_ ), .B2(_04398_ ), .ZN(_01608_ ) );
BUF_X4 _18810_ ( .A(_10578_ ), .Z(_04399_ ) );
NAND4_X1 _18811_ ( .A1(_10668_ ), .A2(_04388_ ), .A3(_04399_ ), .A4(_04382_ ), .ZN(_04400_ ) );
OAI21_X1 _18812_ ( .A(\u_lsu.pmem[2469] ), .B1(_11501_ ), .B2(_04312_ ), .ZN(_04401_ ) );
AOI21_X1 _18813_ ( .A(fanout_net_56 ), .B1(_04400_ ), .B2(_04401_ ), .ZN(_01609_ ) );
OAI21_X1 _18814_ ( .A(\u_lsu.pmem[4196] ), .B1(_03705_ ), .B2(_09919_ ), .ZN(_04402_ ) );
NAND4_X1 _18815_ ( .A1(_09931_ ), .A2(_04376_ ), .A3(_04279_ ), .A4(_02323_ ), .ZN(_04403_ ) );
AOI21_X1 _18816_ ( .A(fanout_net_56 ), .B1(_04402_ ), .B2(_04403_ ), .ZN(_01610_ ) );
NAND4_X1 _18817_ ( .A1(_10671_ ), .A2(_04388_ ), .A3(_04399_ ), .A4(_04382_ ), .ZN(_04404_ ) );
OAI21_X1 _18818_ ( .A(\u_lsu.pmem[2468] ), .B1(_11501_ ), .B2(_04312_ ), .ZN(_04405_ ) );
AOI21_X1 _18819_ ( .A(fanout_net_56 ), .B1(_04404_ ), .B2(_04405_ ), .ZN(_01611_ ) );
NAND4_X1 _18820_ ( .A1(_10674_ ), .A2(_04388_ ), .A3(_04399_ ), .A4(_04382_ ), .ZN(_04406_ ) );
OAI21_X1 _18821_ ( .A(\u_lsu.pmem[2467] ), .B1(_11501_ ), .B2(_04312_ ), .ZN(_04407_ ) );
AOI21_X1 _18822_ ( .A(fanout_net_56 ), .B1(_04406_ ), .B2(_04407_ ), .ZN(_01612_ ) );
BUF_X4 _18823_ ( .A(_04154_ ), .Z(_04408_ ) );
NAND4_X1 _18824_ ( .A1(_10679_ ), .A2(_04388_ ), .A3(_04399_ ), .A4(_04408_ ), .ZN(_04409_ ) );
BUF_X4 _18825_ ( .A(_04265_ ), .Z(_04410_ ) );
OAI21_X1 _18826_ ( .A(\u_lsu.pmem[2466] ), .B1(_11501_ ), .B2(_04410_ ), .ZN(_04411_ ) );
AOI21_X1 _18827_ ( .A(fanout_net_56 ), .B1(_04409_ ), .B2(_04411_ ), .ZN(_01613_ ) );
NAND4_X1 _18828_ ( .A1(_10682_ ), .A2(_04388_ ), .A3(_04399_ ), .A4(_04408_ ), .ZN(_04412_ ) );
OAI21_X1 _18829_ ( .A(\u_lsu.pmem[2465] ), .B1(_11501_ ), .B2(_04410_ ), .ZN(_04413_ ) );
AOI21_X1 _18830_ ( .A(fanout_net_56 ), .B1(_04412_ ), .B2(_04413_ ), .ZN(_01614_ ) );
NAND4_X1 _18831_ ( .A1(_04296_ ), .A2(_10066_ ), .A3(_03753_ ), .A4(_11499_ ), .ZN(_04414_ ) );
OAI21_X1 _18832_ ( .A(\u_lsu.pmem[2464] ), .B1(_11501_ ), .B2(_04410_ ), .ZN(_04415_ ) );
AOI21_X1 _18833_ ( .A(fanout_net_56 ), .B1(_04414_ ), .B2(_04415_ ), .ZN(_01615_ ) );
OAI21_X1 _18834_ ( .A(\u_lsu.pmem[2439] ), .B1(_11521_ ), .B2(_04163_ ), .ZN(_04416_ ) );
NAND4_X1 _18835_ ( .A1(_11542_ ), .A2(_03478_ ), .A3(_04093_ ), .A4(_04094_ ), .ZN(_04417_ ) );
AOI21_X1 _18836_ ( .A(fanout_net_56 ), .B1(_04416_ ), .B2(_04417_ ), .ZN(_01616_ ) );
BUF_X4 _18837_ ( .A(_09647_ ), .Z(_04418_ ) );
OAI21_X1 _18838_ ( .A(\u_lsu.pmem[2438] ), .B1(_11521_ ), .B2(_04418_ ), .ZN(_04419_ ) );
NAND4_X1 _18839_ ( .A1(_11542_ ), .A2(_03056_ ), .A3(_04093_ ), .A4(_04094_ ), .ZN(_04420_ ) );
AOI21_X1 _18840_ ( .A(fanout_net_56 ), .B1(_04419_ ), .B2(_04420_ ), .ZN(_01617_ ) );
OAI21_X1 _18841_ ( .A(\u_lsu.pmem[2437] ), .B1(_11520_ ), .B2(_04418_ ), .ZN(_04421_ ) );
BUF_X4 _18842_ ( .A(_11381_ ), .Z(_04422_ ) );
BUF_X4 _18843_ ( .A(_09522_ ), .Z(_04423_ ) );
NAND4_X1 _18844_ ( .A1(_09512_ ), .A2(_03059_ ), .A3(_04422_ ), .A4(_04423_ ), .ZN(_04424_ ) );
AOI21_X1 _18845_ ( .A(fanout_net_56 ), .B1(_04421_ ), .B2(_04424_ ), .ZN(_01618_ ) );
OAI21_X1 _18846_ ( .A(\u_lsu.pmem[2436] ), .B1(_11520_ ), .B2(_04418_ ), .ZN(_04425_ ) );
NAND4_X1 _18847_ ( .A1(_09512_ ), .A2(_03064_ ), .A3(_04422_ ), .A4(_04423_ ), .ZN(_04426_ ) );
AOI21_X1 _18848_ ( .A(fanout_net_56 ), .B1(_04425_ ), .B2(_04426_ ), .ZN(_01619_ ) );
OAI21_X1 _18849_ ( .A(\u_lsu.pmem[2435] ), .B1(_11520_ ), .B2(_04418_ ), .ZN(_04427_ ) );
NAND4_X1 _18850_ ( .A1(_09512_ ), .A2(_09519_ ), .A3(_04422_ ), .A4(_04423_ ), .ZN(_04428_ ) );
AOI21_X1 _18851_ ( .A(fanout_net_56 ), .B1(_04427_ ), .B2(_04428_ ), .ZN(_01620_ ) );
OAI21_X1 _18852_ ( .A(\u_lsu.pmem[4195] ), .B1(_03705_ ), .B2(_09919_ ), .ZN(_04429_ ) );
NAND4_X1 _18853_ ( .A1(_03091_ ), .A2(_04376_ ), .A3(_04279_ ), .A4(_09916_ ), .ZN(_04430_ ) );
AOI21_X1 _18854_ ( .A(fanout_net_56 ), .B1(_04429_ ), .B2(_04430_ ), .ZN(_01621_ ) );
OAI21_X1 _18855_ ( .A(\u_lsu.pmem[2434] ), .B1(_11520_ ), .B2(_04418_ ), .ZN(_04431_ ) );
NAND4_X1 _18856_ ( .A1(_09537_ ), .A2(_03361_ ), .A3(_04422_ ), .A4(_04423_ ), .ZN(_04432_ ) );
AOI21_X1 _18857_ ( .A(fanout_net_56 ), .B1(_04431_ ), .B2(_04432_ ), .ZN(_01622_ ) );
OAI21_X1 _18858_ ( .A(\u_lsu.pmem[2433] ), .B1(_11520_ ), .B2(_04418_ ), .ZN(_04433_ ) );
NAND4_X1 _18859_ ( .A1(_09512_ ), .A2(_09543_ ), .A3(_04422_ ), .A4(_04423_ ), .ZN(_04434_ ) );
AOI21_X1 _18860_ ( .A(fanout_net_56 ), .B1(_04433_ ), .B2(_04434_ ), .ZN(_01623_ ) );
OAI21_X1 _18861_ ( .A(\u_lsu.pmem[2432] ), .B1(_11520_ ), .B2(_04418_ ), .ZN(_04435_ ) );
NAND4_X1 _18862_ ( .A1(_09512_ ), .A2(_09547_ ), .A3(_04422_ ), .A4(_04423_ ), .ZN(_04436_ ) );
AOI21_X1 _18863_ ( .A(fanout_net_56 ), .B1(_04435_ ), .B2(_04436_ ), .ZN(_01624_ ) );
OAI21_X1 _18864_ ( .A(\u_lsu.pmem[2407] ), .B1(_11547_ ), .B2(_04418_ ), .ZN(_04437_ ) );
NAND3_X1 _18865_ ( .A1(_04161_ ), .A2(_11000_ ), .A3(_11549_ ), .ZN(_04438_ ) );
AOI21_X1 _18866_ ( .A(fanout_net_56 ), .B1(_04437_ ), .B2(_04438_ ), .ZN(_01625_ ) );
OAI21_X1 _18867_ ( .A(\u_lsu.pmem[2406] ), .B1(_11547_ ), .B2(_04418_ ), .ZN(_04439_ ) );
NAND3_X1 _18868_ ( .A1(_04161_ ), .A2(_09579_ ), .A3(_11549_ ), .ZN(_04440_ ) );
AOI21_X1 _18869_ ( .A(fanout_net_56 ), .B1(_04439_ ), .B2(_04440_ ), .ZN(_01626_ ) );
OAI21_X1 _18870_ ( .A(\u_lsu.pmem[2405] ), .B1(_11547_ ), .B2(_04418_ ), .ZN(_04441_ ) );
BUF_X4 _18871_ ( .A(_09641_ ), .Z(_04442_ ) );
NAND3_X1 _18872_ ( .A1(_04442_ ), .A2(_09586_ ), .A3(_11545_ ), .ZN(_04443_ ) );
AOI21_X1 _18873_ ( .A(fanout_net_56 ), .B1(_04441_ ), .B2(_04443_ ), .ZN(_01627_ ) );
BUF_X4 _18874_ ( .A(_09647_ ), .Z(_04444_ ) );
OAI21_X1 _18875_ ( .A(\u_lsu.pmem[2404] ), .B1(_11547_ ), .B2(_04444_ ), .ZN(_04445_ ) );
NAND3_X1 _18876_ ( .A1(_04442_ ), .A2(_09589_ ), .A3(_11545_ ), .ZN(_04446_ ) );
AOI21_X1 _18877_ ( .A(fanout_net_56 ), .B1(_04445_ ), .B2(_04446_ ), .ZN(_01628_ ) );
OAI21_X1 _18878_ ( .A(\u_lsu.pmem[2403] ), .B1(_11547_ ), .B2(_04444_ ), .ZN(_04447_ ) );
NAND3_X1 _18879_ ( .A1(_04442_ ), .A2(_09592_ ), .A3(_11545_ ), .ZN(_04448_ ) );
AOI21_X1 _18880_ ( .A(fanout_net_56 ), .B1(_04447_ ), .B2(_04448_ ), .ZN(_01629_ ) );
OAI21_X1 _18881_ ( .A(\u_lsu.pmem[2402] ), .B1(_11547_ ), .B2(_04444_ ), .ZN(_04449_ ) );
NAND3_X1 _18882_ ( .A1(_04442_ ), .A2(_09695_ ), .A3(_11545_ ), .ZN(_04450_ ) );
AOI21_X1 _18883_ ( .A(fanout_net_56 ), .B1(_04449_ ), .B2(_04450_ ), .ZN(_01630_ ) );
OAI21_X1 _18884_ ( .A(\u_lsu.pmem[2401] ), .B1(_11547_ ), .B2(_04444_ ), .ZN(_04451_ ) );
NAND3_X1 _18885_ ( .A1(_04442_ ), .A2(_09617_ ), .A3(_11545_ ), .ZN(_04452_ ) );
AOI21_X1 _18886_ ( .A(fanout_net_56 ), .B1(_04451_ ), .B2(_04452_ ), .ZN(_01631_ ) );
BUF_X4 _18887_ ( .A(_04210_ ), .Z(_04453_ ) );
BUF_X4 _18888_ ( .A(_03326_ ), .Z(_04454_ ) );
NAND4_X1 _18889_ ( .A1(_09708_ ), .A2(_04453_ ), .A3(_04454_ ), .A4(_04097_ ), .ZN(_04455_ ) );
OAI21_X1 _18890_ ( .A(\u_lsu.pmem[4359] ), .B1(_04071_ ), .B2(_09468_ ), .ZN(_04456_ ) );
AOI21_X1 _18891_ ( .A(fanout_net_56 ), .B1(_04455_ ), .B2(_04456_ ), .ZN(_01632_ ) );
OAI21_X1 _18892_ ( .A(\u_lsu.pmem[4194] ), .B1(_03705_ ), .B2(_09919_ ), .ZN(_04457_ ) );
NAND4_X1 _18893_ ( .A1(_09938_ ), .A2(_04376_ ), .A3(_04279_ ), .A4(_09916_ ), .ZN(_04458_ ) );
AOI21_X1 _18894_ ( .A(fanout_net_56 ), .B1(_04457_ ), .B2(_04458_ ), .ZN(_01633_ ) );
OAI21_X1 _18895_ ( .A(\u_lsu.pmem[2400] ), .B1(_11547_ ), .B2(_04444_ ), .ZN(_04459_ ) );
NAND3_X1 _18896_ ( .A1(_04442_ ), .A2(_09622_ ), .A3(_11545_ ), .ZN(_04460_ ) );
AOI21_X1 _18897_ ( .A(fanout_net_56 ), .B1(_04459_ ), .B2(_04460_ ), .ZN(_01634_ ) );
OAI21_X1 _18898_ ( .A(\u_lsu.pmem[2375] ), .B1(_11572_ ), .B2(_04444_ ), .ZN(_04461_ ) );
NAND3_X1 _18899_ ( .A1(_04442_ ), .A2(_10330_ ), .A3(_11574_ ), .ZN(_04462_ ) );
AOI21_X1 _18900_ ( .A(fanout_net_56 ), .B1(_04461_ ), .B2(_04462_ ), .ZN(_01635_ ) );
OAI21_X1 _18901_ ( .A(\u_lsu.pmem[2374] ), .B1(_11572_ ), .B2(_04444_ ), .ZN(_04463_ ) );
NAND3_X1 _18902_ ( .A1(_04442_ ), .A2(_09579_ ), .A3(_11574_ ), .ZN(_04464_ ) );
AOI21_X1 _18903_ ( .A(fanout_net_56 ), .B1(_04463_ ), .B2(_04464_ ), .ZN(_01636_ ) );
OAI21_X1 _18904_ ( .A(\u_lsu.pmem[2373] ), .B1(_11572_ ), .B2(_04444_ ), .ZN(_04465_ ) );
NAND3_X1 _18905_ ( .A1(_04442_ ), .A2(_09586_ ), .A3(_11570_ ), .ZN(_04466_ ) );
AOI21_X1 _18906_ ( .A(fanout_net_56 ), .B1(_04465_ ), .B2(_04466_ ), .ZN(_01637_ ) );
OAI21_X1 _18907_ ( .A(\u_lsu.pmem[2372] ), .B1(_11572_ ), .B2(_04444_ ), .ZN(_04467_ ) );
NAND3_X1 _18908_ ( .A1(_04442_ ), .A2(_10486_ ), .A3(_11570_ ), .ZN(_04468_ ) );
AOI21_X1 _18909_ ( .A(fanout_net_57 ), .B1(_04467_ ), .B2(_04468_ ), .ZN(_01638_ ) );
OAI21_X1 _18910_ ( .A(\u_lsu.pmem[2371] ), .B1(_11572_ ), .B2(_04444_ ), .ZN(_04469_ ) );
BUF_X4 _18911_ ( .A(_09641_ ), .Z(_04470_ ) );
NAND3_X1 _18912_ ( .A1(_04470_ ), .A2(_09592_ ), .A3(_11570_ ), .ZN(_04471_ ) );
AOI21_X1 _18913_ ( .A(fanout_net_57 ), .B1(_04469_ ), .B2(_04471_ ), .ZN(_01639_ ) );
BUF_X4 _18914_ ( .A(_10720_ ), .Z(_04472_ ) );
OAI21_X1 _18915_ ( .A(\u_lsu.pmem[2370] ), .B1(_11572_ ), .B2(_04472_ ), .ZN(_04473_ ) );
NAND3_X1 _18916_ ( .A1(_04470_ ), .A2(_09695_ ), .A3(_11570_ ), .ZN(_04474_ ) );
AOI21_X1 _18917_ ( .A(fanout_net_57 ), .B1(_04473_ ), .B2(_04474_ ), .ZN(_01640_ ) );
OAI21_X1 _18918_ ( .A(\u_lsu.pmem[2369] ), .B1(_11572_ ), .B2(_04472_ ), .ZN(_04475_ ) );
NAND3_X1 _18919_ ( .A1(_04470_ ), .A2(_09617_ ), .A3(_11570_ ), .ZN(_04476_ ) );
AOI21_X1 _18920_ ( .A(fanout_net_57 ), .B1(_04475_ ), .B2(_04476_ ), .ZN(_01641_ ) );
OAI21_X1 _18921_ ( .A(\u_lsu.pmem[2368] ), .B1(_11572_ ), .B2(_04472_ ), .ZN(_04477_ ) );
NAND3_X1 _18922_ ( .A1(_04470_ ), .A2(_09622_ ), .A3(_11570_ ), .ZN(_04478_ ) );
AOI21_X1 _18923_ ( .A(fanout_net_57 ), .B1(_04477_ ), .B2(_04478_ ), .ZN(_01642_ ) );
NAND4_X1 _18924_ ( .A1(_09670_ ), .A2(_04453_ ), .A3(_04399_ ), .A4(_04408_ ), .ZN(_04479_ ) );
OAI21_X1 _18925_ ( .A(\u_lsu.pmem[2343] ), .B1(_11597_ ), .B2(_04410_ ), .ZN(_04480_ ) );
AOI21_X1 _18926_ ( .A(fanout_net_57 ), .B1(_04479_ ), .B2(_04480_ ), .ZN(_01643_ ) );
OAI21_X1 _18927_ ( .A(\u_lsu.pmem[4193] ), .B1(_03705_ ), .B2(_09919_ ), .ZN(_04481_ ) );
NAND4_X1 _18928_ ( .A1(_03143_ ), .A2(_04376_ ), .A3(_04279_ ), .A4(_09916_ ), .ZN(_04482_ ) );
AOI21_X1 _18929_ ( .A(fanout_net_57 ), .B1(_04481_ ), .B2(_04482_ ), .ZN(_01644_ ) );
NAND4_X1 _18930_ ( .A1(_09681_ ), .A2(_04453_ ), .A3(_04399_ ), .A4(_04408_ ), .ZN(_04483_ ) );
OAI21_X1 _18931_ ( .A(\u_lsu.pmem[2342] ), .B1(_11597_ ), .B2(_04410_ ), .ZN(_04484_ ) );
AOI21_X1 _18932_ ( .A(fanout_net_57 ), .B1(_04483_ ), .B2(_04484_ ), .ZN(_01645_ ) );
NAND4_X1 _18933_ ( .A1(_09685_ ), .A2(_04453_ ), .A3(_04399_ ), .A4(_04408_ ), .ZN(_04485_ ) );
OAI21_X1 _18934_ ( .A(\u_lsu.pmem[2341] ), .B1(_11597_ ), .B2(_04410_ ), .ZN(_04486_ ) );
AOI21_X1 _18935_ ( .A(fanout_net_57 ), .B1(_04485_ ), .B2(_04486_ ), .ZN(_01646_ ) );
NOR2_X4 _18936_ ( .A1(_11597_ ), .A2(_09635_ ), .ZN(_04487_ ) );
OAI21_X1 _18937_ ( .A(_09109_ ), .B1(_04487_ ), .B2(\u_lsu.pmem[2340] ), .ZN(_04488_ ) );
AOI21_X1 _18938_ ( .A(_04488_ ), .B1(_09149_ ), .B2(_04487_ ), .ZN(_01647_ ) );
OAI21_X1 _18939_ ( .A(\u_lsu.pmem[2339] ), .B1(_11598_ ), .B2(_04472_ ), .ZN(_04489_ ) );
NAND3_X1 _18940_ ( .A1(_04470_ ), .A2(_09592_ ), .A3(_11596_ ), .ZN(_04490_ ) );
AOI21_X1 _18941_ ( .A(fanout_net_57 ), .B1(_04489_ ), .B2(_04490_ ), .ZN(_01648_ ) );
OAI21_X1 _18942_ ( .A(\u_lsu.pmem[2338] ), .B1(_11598_ ), .B2(_04472_ ), .ZN(_04491_ ) );
NAND3_X1 _18943_ ( .A1(_04470_ ), .A2(_09695_ ), .A3(_11596_ ), .ZN(_04492_ ) );
AOI21_X1 _18944_ ( .A(fanout_net_57 ), .B1(_04491_ ), .B2(_04492_ ), .ZN(_01649_ ) );
OAI21_X1 _18945_ ( .A(\u_lsu.pmem[2337] ), .B1(_11598_ ), .B2(_04472_ ), .ZN(_04493_ ) );
NAND3_X1 _18946_ ( .A1(_04470_ ), .A2(_09617_ ), .A3(_11596_ ), .ZN(_04494_ ) );
AOI21_X1 _18947_ ( .A(fanout_net_57 ), .B1(_04493_ ), .B2(_04494_ ), .ZN(_01650_ ) );
NAND4_X1 _18948_ ( .A1(_09703_ ), .A2(_04453_ ), .A3(_04399_ ), .A4(_04408_ ), .ZN(_04495_ ) );
OAI21_X1 _18949_ ( .A(\u_lsu.pmem[2336] ), .B1(_11597_ ), .B2(_04410_ ), .ZN(_04496_ ) );
AOI21_X1 _18950_ ( .A(fanout_net_57 ), .B1(_04495_ ), .B2(_04496_ ), .ZN(_01651_ ) );
NAND4_X1 _18951_ ( .A1(_09708_ ), .A2(_04453_ ), .A3(_04399_ ), .A4(_04408_ ), .ZN(_04497_ ) );
OAI21_X1 _18952_ ( .A(\u_lsu.pmem[2311] ), .B1(_04386_ ), .B2(_02200_ ), .ZN(_04498_ ) );
AOI21_X1 _18953_ ( .A(fanout_net_57 ), .B1(_04497_ ), .B2(_04498_ ), .ZN(_01652_ ) );
BUF_X4 _18954_ ( .A(_10578_ ), .Z(_04499_ ) );
NAND4_X1 _18955_ ( .A1(_09715_ ), .A2(_04453_ ), .A3(_04499_ ), .A4(_04408_ ), .ZN(_04500_ ) );
OAI21_X1 _18956_ ( .A(\u_lsu.pmem[2310] ), .B1(_04386_ ), .B2(_02200_ ), .ZN(_04501_ ) );
AOI21_X1 _18957_ ( .A(fanout_net_57 ), .B1(_04500_ ), .B2(_04501_ ), .ZN(_01653_ ) );
NAND4_X1 _18958_ ( .A1(_09718_ ), .A2(_04453_ ), .A3(_04499_ ), .A4(_04408_ ), .ZN(_04502_ ) );
OAI21_X1 _18959_ ( .A(\u_lsu.pmem[2309] ), .B1(_04386_ ), .B2(_02199_ ), .ZN(_04503_ ) );
AOI21_X1 _18960_ ( .A(fanout_net_57 ), .B1(_04502_ ), .B2(_04503_ ), .ZN(_01654_ ) );
OAI21_X1 _18961_ ( .A(\u_lsu.pmem[4192] ), .B1(_03705_ ), .B2(_09919_ ), .ZN(_04504_ ) );
NAND4_X1 _18962_ ( .A1(_09944_ ), .A2(_04376_ ), .A3(_04279_ ), .A4(_09916_ ), .ZN(_04505_ ) );
AOI21_X1 _18963_ ( .A(fanout_net_57 ), .B1(_04504_ ), .B2(_04505_ ), .ZN(_01655_ ) );
NAND4_X1 _18964_ ( .A1(_09721_ ), .A2(_04453_ ), .A3(_04499_ ), .A4(_04408_ ), .ZN(_04506_ ) );
OAI21_X1 _18965_ ( .A(\u_lsu.pmem[2308] ), .B1(_04386_ ), .B2(_02199_ ), .ZN(_04507_ ) );
AOI21_X1 _18966_ ( .A(fanout_net_57 ), .B1(_04506_ ), .B2(_04507_ ), .ZN(_01656_ ) );
BUF_X4 _18967_ ( .A(_04154_ ), .Z(_04508_ ) );
NAND4_X1 _18968_ ( .A1(_09725_ ), .A2(_04453_ ), .A3(_04499_ ), .A4(_04508_ ), .ZN(_04509_ ) );
OAI21_X1 _18969_ ( .A(\u_lsu.pmem[2307] ), .B1(_04386_ ), .B2(_02199_ ), .ZN(_04510_ ) );
AOI21_X1 _18970_ ( .A(fanout_net_57 ), .B1(_04509_ ), .B2(_04510_ ), .ZN(_01657_ ) );
OR3_X2 _18971_ ( .A1(_11159_ ), .A2(_02199_ ), .A3(_09973_ ), .ZN(_04511_ ) );
OAI21_X1 _18972_ ( .A(\u_lsu.pmem[2306] ), .B1(_04386_ ), .B2(_02199_ ), .ZN(_04512_ ) );
AOI21_X1 _18973_ ( .A(fanout_net_57 ), .B1(_04511_ ), .B2(_04512_ ), .ZN(_01658_ ) );
BUF_X4 _18974_ ( .A(_04210_ ), .Z(_04513_ ) );
NAND4_X1 _18975_ ( .A1(_09733_ ), .A2(_04513_ ), .A3(_04499_ ), .A4(_04508_ ), .ZN(_04514_ ) );
BUF_X4 _18976_ ( .A(_03919_ ), .Z(_04515_ ) );
OAI21_X1 _18977_ ( .A(\u_lsu.pmem[2305] ), .B1(_04515_ ), .B2(_02199_ ), .ZN(_04516_ ) );
AOI21_X1 _18978_ ( .A(fanout_net_57 ), .B1(_04514_ ), .B2(_04516_ ), .ZN(_01659_ ) );
NAND4_X1 _18979_ ( .A1(_09736_ ), .A2(_04513_ ), .A3(_04499_ ), .A4(_04508_ ), .ZN(_04517_ ) );
OAI21_X1 _18980_ ( .A(\u_lsu.pmem[2304] ), .B1(_04515_ ), .B2(_02199_ ), .ZN(_04518_ ) );
AOI21_X1 _18981_ ( .A(fanout_net_57 ), .B1(_04517_ ), .B2(_04518_ ), .ZN(_01660_ ) );
NOR2_X1 _18982_ ( .A1(_03850_ ), .A2(_02221_ ), .ZN(_04519_ ) );
NOR2_X1 _18983_ ( .A1(_04519_ ), .A2(\u_lsu.pmem[2279] ), .ZN(_04520_ ) );
AOI211_X1 _18984_ ( .A(fanout_net_57 ), .B(_04520_ ), .C1(_04216_ ), .C2(_04519_ ), .ZN(_01661_ ) );
NAND4_X1 _18985_ ( .A1(_09756_ ), .A2(_04513_ ), .A3(_04499_ ), .A4(_04508_ ), .ZN(_04521_ ) );
OAI21_X1 _18986_ ( .A(\u_lsu.pmem[2278] ), .B1(_04515_ ), .B2(_02222_ ), .ZN(_04522_ ) );
AOI21_X1 _18987_ ( .A(fanout_net_57 ), .B1(_04521_ ), .B2(_04522_ ), .ZN(_01662_ ) );
NAND4_X1 _18988_ ( .A1(_09763_ ), .A2(_04513_ ), .A3(_04499_ ), .A4(_04508_ ), .ZN(_04523_ ) );
OAI21_X1 _18989_ ( .A(\u_lsu.pmem[2277] ), .B1(_04515_ ), .B2(_02222_ ), .ZN(_04524_ ) );
AOI21_X1 _18990_ ( .A(fanout_net_57 ), .B1(_04523_ ), .B2(_04524_ ), .ZN(_01663_ ) );
NAND4_X1 _18991_ ( .A1(_09770_ ), .A2(_04513_ ), .A3(_04499_ ), .A4(_04508_ ), .ZN(_04525_ ) );
OAI21_X1 _18992_ ( .A(\u_lsu.pmem[2276] ), .B1(_04515_ ), .B2(_02221_ ), .ZN(_04526_ ) );
AOI21_X1 _18993_ ( .A(fanout_net_57 ), .B1(_04525_ ), .B2(_04526_ ), .ZN(_01664_ ) );
NAND4_X1 _18994_ ( .A1(_09775_ ), .A2(_04513_ ), .A3(_04499_ ), .A4(_04508_ ), .ZN(_04527_ ) );
OAI21_X1 _18995_ ( .A(\u_lsu.pmem[2275] ), .B1(_04515_ ), .B2(_02221_ ), .ZN(_04528_ ) );
AOI21_X1 _18996_ ( .A(fanout_net_57 ), .B1(_04527_ ), .B2(_04528_ ), .ZN(_01665_ ) );
OR3_X1 _18997_ ( .A1(_09567_ ), .A2(_09459_ ), .A3(_09949_ ), .ZN(_04529_ ) );
OAI21_X1 _18998_ ( .A(\u_lsu.pmem[4167] ), .B1(_04071_ ), .B2(_09949_ ), .ZN(_04530_ ) );
AOI21_X1 _18999_ ( .A(fanout_net_57 ), .B1(_04529_ ), .B2(_04530_ ), .ZN(_01666_ ) );
BUF_X4 _19000_ ( .A(_10578_ ), .Z(_04531_ ) );
NAND4_X1 _19001_ ( .A1(_09780_ ), .A2(_04513_ ), .A3(_04531_ ), .A4(_04508_ ), .ZN(_04532_ ) );
OAI21_X1 _19002_ ( .A(\u_lsu.pmem[2274] ), .B1(_04515_ ), .B2(_02221_ ), .ZN(_04533_ ) );
AOI21_X1 _19003_ ( .A(fanout_net_57 ), .B1(_04532_ ), .B2(_04533_ ), .ZN(_01667_ ) );
NAND4_X1 _19004_ ( .A1(_09787_ ), .A2(_04513_ ), .A3(_04531_ ), .A4(_04508_ ), .ZN(_04534_ ) );
OAI21_X1 _19005_ ( .A(\u_lsu.pmem[2273] ), .B1(_04515_ ), .B2(_02221_ ), .ZN(_04535_ ) );
AOI21_X1 _19006_ ( .A(fanout_net_57 ), .B1(_04534_ ), .B2(_04535_ ), .ZN(_01668_ ) );
NAND4_X1 _19007_ ( .A1(_09791_ ), .A2(_04513_ ), .A3(_04531_ ), .A4(_04508_ ), .ZN(_04536_ ) );
OAI21_X1 _19008_ ( .A(\u_lsu.pmem[2272] ), .B1(_04515_ ), .B2(_02221_ ), .ZN(_04537_ ) );
AOI21_X1 _19009_ ( .A(fanout_net_58 ), .B1(_04536_ ), .B2(_04537_ ), .ZN(_01669_ ) );
NOR2_X1 _19010_ ( .A1(_03850_ ), .A2(_02243_ ), .ZN(_04538_ ) );
NOR2_X1 _19011_ ( .A1(_04538_ ), .A2(\u_lsu.pmem[2247] ), .ZN(_04539_ ) );
AOI211_X1 _19012_ ( .A(fanout_net_58 ), .B(_04539_ ), .C1(_04216_ ), .C2(_04538_ ), .ZN(_01670_ ) );
BUF_X4 _19013_ ( .A(_04154_ ), .Z(_04540_ ) );
NAND4_X1 _19014_ ( .A1(_09804_ ), .A2(_09806_ ), .A3(_04531_ ), .A4(_04540_ ), .ZN(_04541_ ) );
OAI21_X1 _19015_ ( .A(\u_lsu.pmem[2246] ), .B1(_04515_ ), .B2(_02244_ ), .ZN(_04542_ ) );
AOI21_X1 _19016_ ( .A(fanout_net_58 ), .B1(_04541_ ), .B2(_04542_ ), .ZN(_01671_ ) );
NAND4_X1 _19017_ ( .A1(_09811_ ), .A2(_04513_ ), .A3(_04531_ ), .A4(_04540_ ), .ZN(_04543_ ) );
BUF_X4 _19018_ ( .A(_03919_ ), .Z(_04544_ ) );
OAI21_X1 _19019_ ( .A(\u_lsu.pmem[2245] ), .B1(_04544_ ), .B2(_02244_ ), .ZN(_04545_ ) );
AOI21_X1 _19020_ ( .A(fanout_net_58 ), .B1(_04543_ ), .B2(_04545_ ), .ZN(_01672_ ) );
BUF_X4 _19021_ ( .A(_04210_ ), .Z(_04546_ ) );
NAND4_X1 _19022_ ( .A1(_09815_ ), .A2(_04546_ ), .A3(_04531_ ), .A4(_04540_ ), .ZN(_04547_ ) );
OAI21_X1 _19023_ ( .A(\u_lsu.pmem[2244] ), .B1(_04544_ ), .B2(_02243_ ), .ZN(_04548_ ) );
AOI21_X1 _19024_ ( .A(fanout_net_58 ), .B1(_04547_ ), .B2(_04548_ ), .ZN(_01673_ ) );
NAND4_X1 _19025_ ( .A1(_09819_ ), .A2(_04546_ ), .A3(_04531_ ), .A4(_04540_ ), .ZN(_04549_ ) );
OAI21_X1 _19026_ ( .A(\u_lsu.pmem[2243] ), .B1(_04544_ ), .B2(_02243_ ), .ZN(_04550_ ) );
AOI21_X1 _19027_ ( .A(fanout_net_58 ), .B1(_04549_ ), .B2(_04550_ ), .ZN(_01674_ ) );
NAND4_X1 _19028_ ( .A1(_09827_ ), .A2(_04546_ ), .A3(_04531_ ), .A4(_04540_ ), .ZN(_04551_ ) );
OAI21_X1 _19029_ ( .A(\u_lsu.pmem[2242] ), .B1(_04544_ ), .B2(_02243_ ), .ZN(_04552_ ) );
AOI21_X1 _19030_ ( .A(fanout_net_58 ), .B1(_04551_ ), .B2(_04552_ ), .ZN(_01675_ ) );
NAND4_X1 _19031_ ( .A1(_09831_ ), .A2(_04546_ ), .A3(_04531_ ), .A4(_04540_ ), .ZN(_04553_ ) );
OAI21_X1 _19032_ ( .A(\u_lsu.pmem[2241] ), .B1(_04544_ ), .B2(_02243_ ), .ZN(_04554_ ) );
AOI21_X1 _19033_ ( .A(fanout_net_58 ), .B1(_04553_ ), .B2(_04554_ ), .ZN(_01676_ ) );
OAI21_X1 _19034_ ( .A(\u_lsu.pmem[4166] ), .B1(_03705_ ), .B2(_09959_ ), .ZN(_04555_ ) );
BUF_X4 _19035_ ( .A(_09455_ ), .Z(_04556_ ) );
NAND4_X1 _19036_ ( .A1(_09957_ ), .A2(_03361_ ), .A3(_04556_ ), .A4(_03646_ ), .ZN(_04557_ ) );
AOI21_X1 _19037_ ( .A(fanout_net_58 ), .B1(_04555_ ), .B2(_04557_ ), .ZN(_01677_ ) );
NAND4_X1 _19038_ ( .A1(_09835_ ), .A2(_04546_ ), .A3(_04531_ ), .A4(_04540_ ), .ZN(_04558_ ) );
OAI21_X1 _19039_ ( .A(\u_lsu.pmem[2240] ), .B1(_04544_ ), .B2(_02243_ ), .ZN(_04559_ ) );
AOI21_X1 _19040_ ( .A(fanout_net_58 ), .B1(_04558_ ), .B2(_04559_ ), .ZN(_01678_ ) );
BUF_X4 _19041_ ( .A(_10578_ ), .Z(_04560_ ) );
NAND4_X1 _19042_ ( .A1(_09840_ ), .A2(_04546_ ), .A3(_04560_ ), .A4(_04540_ ), .ZN(_04561_ ) );
OAI21_X1 _19043_ ( .A(\u_lsu.pmem[2215] ), .B1(_04544_ ), .B2(_02270_ ), .ZN(_04562_ ) );
AOI21_X1 _19044_ ( .A(fanout_net_58 ), .B1(_04561_ ), .B2(_04562_ ), .ZN(_01679_ ) );
NAND4_X1 _19045_ ( .A1(_09849_ ), .A2(_04546_ ), .A3(_04560_ ), .A4(_04540_ ), .ZN(_04563_ ) );
OAI21_X1 _19046_ ( .A(\u_lsu.pmem[2214] ), .B1(_04544_ ), .B2(_02270_ ), .ZN(_04564_ ) );
AOI21_X1 _19047_ ( .A(fanout_net_58 ), .B1(_04563_ ), .B2(_04564_ ), .ZN(_01680_ ) );
NAND4_X1 _19048_ ( .A1(_09853_ ), .A2(_04546_ ), .A3(_04560_ ), .A4(_04540_ ), .ZN(_04565_ ) );
OAI21_X1 _19049_ ( .A(\u_lsu.pmem[2213] ), .B1(_04544_ ), .B2(_02269_ ), .ZN(_04566_ ) );
AOI21_X1 _19050_ ( .A(fanout_net_58 ), .B1(_04565_ ), .B2(_04566_ ), .ZN(_01681_ ) );
BUF_X4 _19051_ ( .A(_04154_ ), .Z(_04567_ ) );
NAND4_X1 _19052_ ( .A1(_09858_ ), .A2(_04546_ ), .A3(_04560_ ), .A4(_04567_ ), .ZN(_04568_ ) );
OAI21_X1 _19053_ ( .A(\u_lsu.pmem[2212] ), .B1(_04544_ ), .B2(_02269_ ), .ZN(_04569_ ) );
AOI21_X1 _19054_ ( .A(fanout_net_58 ), .B1(_04568_ ), .B2(_04569_ ), .ZN(_01682_ ) );
NAND4_X1 _19055_ ( .A1(_09861_ ), .A2(_04546_ ), .A3(_04560_ ), .A4(_04567_ ), .ZN(_04570_ ) );
BUF_X8 _19056_ ( .A(_09471_ ), .Z(_04571_ ) );
BUF_X4 _19057_ ( .A(_04571_ ), .Z(_04572_ ) );
OAI21_X1 _19058_ ( .A(\u_lsu.pmem[2211] ), .B1(_04572_ ), .B2(_02269_ ), .ZN(_04573_ ) );
AOI21_X1 _19059_ ( .A(fanout_net_58 ), .B1(_04570_ ), .B2(_04573_ ), .ZN(_01683_ ) );
BUF_X4 _19060_ ( .A(_04210_ ), .Z(_04574_ ) );
NAND4_X1 _19061_ ( .A1(_09864_ ), .A2(_04574_ ), .A3(_04560_ ), .A4(_04567_ ), .ZN(_04575_ ) );
OAI21_X1 _19062_ ( .A(\u_lsu.pmem[2210] ), .B1(_04572_ ), .B2(_02269_ ), .ZN(_04576_ ) );
AOI21_X1 _19063_ ( .A(fanout_net_58 ), .B1(_04575_ ), .B2(_04576_ ), .ZN(_01684_ ) );
NAND4_X1 _19064_ ( .A1(_09867_ ), .A2(_04574_ ), .A3(_04560_ ), .A4(_04567_ ), .ZN(_04577_ ) );
OAI21_X1 _19065_ ( .A(\u_lsu.pmem[2209] ), .B1(_04572_ ), .B2(_02269_ ), .ZN(_04578_ ) );
AOI21_X1 _19066_ ( .A(fanout_net_58 ), .B1(_04577_ ), .B2(_04578_ ), .ZN(_01685_ ) );
NAND4_X1 _19067_ ( .A1(_09881_ ), .A2(_09676_ ), .A3(_09979_ ), .A4(_03978_ ), .ZN(_04579_ ) );
OAI21_X1 _19068_ ( .A(\u_lsu.pmem[2208] ), .B1(_04572_ ), .B2(_02269_ ), .ZN(_04580_ ) );
AOI21_X1 _19069_ ( .A(fanout_net_58 ), .B1(_04579_ ), .B2(_04580_ ), .ZN(_01686_ ) );
OAI21_X1 _19070_ ( .A(\u_lsu.pmem[2183] ), .B1(_02293_ ), .B2(_04472_ ), .ZN(_04581_ ) );
NAND4_X1 _19071_ ( .A1(_09893_ ), .A2(_03478_ ), .A3(_04422_ ), .A4(_04423_ ), .ZN(_04582_ ) );
AOI21_X1 _19072_ ( .A(fanout_net_58 ), .B1(_04581_ ), .B2(_04582_ ), .ZN(_01687_ ) );
BUF_X4 _19073_ ( .A(_09459_ ), .Z(_04583_ ) );
OAI21_X1 _19074_ ( .A(\u_lsu.pmem[4165] ), .B1(_04583_ ), .B2(_09959_ ), .ZN(_04584_ ) );
BUF_X4 _19075_ ( .A(_09539_ ), .Z(_04585_ ) );
NAND4_X1 _19076_ ( .A1(_09961_ ), .A2(_04585_ ), .A3(_04556_ ), .A4(_11159_ ), .ZN(_04586_ ) );
AOI21_X1 _19077_ ( .A(fanout_net_58 ), .B1(_04584_ ), .B2(_04586_ ), .ZN(_01688_ ) );
OAI21_X1 _19078_ ( .A(\u_lsu.pmem[2182] ), .B1(_02293_ ), .B2(_04472_ ), .ZN(_04587_ ) );
NAND4_X1 _19079_ ( .A1(_09893_ ), .A2(_03056_ ), .A3(_04422_ ), .A4(_04423_ ), .ZN(_04588_ ) );
AOI21_X1 _19080_ ( .A(fanout_net_58 ), .B1(_04587_ ), .B2(_04588_ ), .ZN(_01689_ ) );
OAI21_X1 _19081_ ( .A(\u_lsu.pmem[2181] ), .B1(_02292_ ), .B2(_04472_ ), .ZN(_04589_ ) );
NAND4_X1 _19082_ ( .A1(_09893_ ), .A2(_03059_ ), .A3(_04422_ ), .A4(_04423_ ), .ZN(_04590_ ) );
AOI21_X1 _19083_ ( .A(fanout_net_58 ), .B1(_04589_ ), .B2(_04590_ ), .ZN(_01690_ ) );
OAI21_X1 _19084_ ( .A(\u_lsu.pmem[2180] ), .B1(_02292_ ), .B2(_04472_ ), .ZN(_04591_ ) );
NAND4_X1 _19085_ ( .A1(_09893_ ), .A2(_03064_ ), .A3(_04422_ ), .A4(_04423_ ), .ZN(_04592_ ) );
AOI21_X1 _19086_ ( .A(fanout_net_58 ), .B1(_04591_ ), .B2(_04592_ ), .ZN(_01691_ ) );
BUF_X4 _19087_ ( .A(_10720_ ), .Z(_04593_ ) );
OAI21_X1 _19088_ ( .A(\u_lsu.pmem[2179] ), .B1(_02292_ ), .B2(_04593_ ), .ZN(_04594_ ) );
BUF_X4 _19089_ ( .A(_09522_ ), .Z(_04595_ ) );
NAND4_X1 _19090_ ( .A1(_09893_ ), .A2(_09519_ ), .A3(_10065_ ), .A4(_04595_ ), .ZN(_04596_ ) );
AOI21_X1 _19091_ ( .A(fanout_net_58 ), .B1(_04594_ ), .B2(_04596_ ), .ZN(_01692_ ) );
OAI21_X1 _19092_ ( .A(\u_lsu.pmem[2178] ), .B1(_02292_ ), .B2(_04593_ ), .ZN(_04597_ ) );
NAND4_X1 _19093_ ( .A1(_09906_ ), .A2(_04585_ ), .A3(_10065_ ), .A4(_04595_ ), .ZN(_04598_ ) );
AOI21_X1 _19094_ ( .A(fanout_net_58 ), .B1(_04597_ ), .B2(_04598_ ), .ZN(_01693_ ) );
OAI21_X1 _19095_ ( .A(\u_lsu.pmem[2177] ), .B1(_02292_ ), .B2(_04593_ ), .ZN(_04599_ ) );
NAND4_X1 _19096_ ( .A1(_09893_ ), .A2(_09543_ ), .A3(_10065_ ), .A4(_04595_ ), .ZN(_04600_ ) );
AOI21_X1 _19097_ ( .A(fanout_net_58 ), .B1(_04599_ ), .B2(_04600_ ), .ZN(_01694_ ) );
OAI21_X1 _19098_ ( .A(\u_lsu.pmem[2176] ), .B1(_02292_ ), .B2(_04593_ ), .ZN(_04601_ ) );
NAND4_X1 _19099_ ( .A1(_09893_ ), .A2(_09547_ ), .A3(_10065_ ), .A4(_04595_ ), .ZN(_04602_ ) );
AOI21_X1 _19100_ ( .A(fanout_net_58 ), .B1(_04601_ ), .B2(_04602_ ), .ZN(_01695_ ) );
NOR2_X4 _19101_ ( .A1(_09450_ ), .A2(_02315_ ), .ZN(_04603_ ) );
NOR2_X1 _19102_ ( .A1(_04603_ ), .A2(\u_lsu.pmem[2151] ), .ZN(_04604_ ) );
AOI211_X1 _19103_ ( .A(fanout_net_58 ), .B(_04604_ ), .C1(_04216_ ), .C2(_04603_ ), .ZN(_01696_ ) );
NAND2_X1 _19104_ ( .A1(_04603_ ), .A2(_11145_ ), .ZN(_04605_ ) );
OAI21_X1 _19105_ ( .A(\u_lsu.pmem[2150] ), .B1(_04572_ ), .B2(_02316_ ), .ZN(_04606_ ) );
AOI21_X1 _19106_ ( .A(fanout_net_58 ), .B1(_04605_ ), .B2(_04606_ ), .ZN(_01697_ ) );
NAND2_X1 _19107_ ( .A1(_04603_ ), .A2(_11148_ ), .ZN(_04607_ ) );
OAI21_X1 _19108_ ( .A(\u_lsu.pmem[2149] ), .B1(_04572_ ), .B2(_02316_ ), .ZN(_04608_ ) );
AOI21_X1 _19109_ ( .A(fanout_net_58 ), .B1(_04607_ ), .B2(_04608_ ), .ZN(_01698_ ) );
OAI21_X1 _19110_ ( .A(\u_lsu.pmem[4164] ), .B1(_04583_ ), .B2(_09959_ ), .ZN(_04609_ ) );
NAND4_X1 _19111_ ( .A1(_09966_ ), .A2(_04585_ ), .A3(_04556_ ), .A4(_11159_ ), .ZN(_04610_ ) );
AOI21_X1 _19112_ ( .A(fanout_net_59 ), .B1(_04609_ ), .B2(_04610_ ), .ZN(_01699_ ) );
NAND2_X1 _19113_ ( .A1(_04603_ ), .A2(_03084_ ), .ZN(_04611_ ) );
OAI21_X1 _19114_ ( .A(\u_lsu.pmem[2148] ), .B1(_04572_ ), .B2(_02315_ ), .ZN(_04612_ ) );
AOI21_X1 _19115_ ( .A(fanout_net_59 ), .B1(_04611_ ), .B2(_04612_ ), .ZN(_01700_ ) );
NAND2_X1 _19116_ ( .A1(_04603_ ), .A2(_03114_ ), .ZN(_04613_ ) );
OAI21_X1 _19117_ ( .A(\u_lsu.pmem[2147] ), .B1(_04572_ ), .B2(_02315_ ), .ZN(_04614_ ) );
AOI21_X1 _19118_ ( .A(fanout_net_59 ), .B1(_04613_ ), .B2(_04614_ ), .ZN(_01701_ ) );
NAND2_X1 _19119_ ( .A1(_04603_ ), .A2(_03145_ ), .ZN(_04615_ ) );
OAI21_X1 _19120_ ( .A(\u_lsu.pmem[2146] ), .B1(_04572_ ), .B2(_02315_ ), .ZN(_04616_ ) );
AOI21_X1 _19121_ ( .A(fanout_net_59 ), .B1(_04615_ ), .B2(_04616_ ), .ZN(_01702_ ) );
NAND2_X1 _19122_ ( .A1(_04603_ ), .A2(_03174_ ), .ZN(_04617_ ) );
OAI21_X1 _19123_ ( .A(\u_lsu.pmem[2145] ), .B1(_04572_ ), .B2(_02315_ ), .ZN(_04618_ ) );
AOI21_X1 _19124_ ( .A(fanout_net_59 ), .B1(_04617_ ), .B2(_04618_ ), .ZN(_01703_ ) );
NAND2_X1 _19125_ ( .A1(_04603_ ), .A2(_03203_ ), .ZN(_04619_ ) );
BUF_X4 _19126_ ( .A(_04571_ ), .Z(_04620_ ) );
OAI21_X1 _19127_ ( .A(\u_lsu.pmem[2144] ), .B1(_04620_ ), .B2(_02315_ ), .ZN(_04621_ ) );
AOI21_X1 _19128_ ( .A(fanout_net_59 ), .B1(_04619_ ), .B2(_04621_ ), .ZN(_01704_ ) );
NOR2_X1 _19129_ ( .A1(_03850_ ), .A2(_02337_ ), .ZN(_04622_ ) );
NOR2_X1 _19130_ ( .A1(_04622_ ), .A2(\u_lsu.pmem[2119] ), .ZN(_04623_ ) );
AOI211_X1 _19131_ ( .A(fanout_net_59 ), .B(_04623_ ), .C1(_04216_ ), .C2(_04622_ ), .ZN(_01705_ ) );
NAND4_X1 _19132_ ( .A1(_04296_ ), .A2(_09957_ ), .A3(_09979_ ), .A4(_03978_ ), .ZN(_04624_ ) );
OAI21_X1 _19133_ ( .A(\u_lsu.pmem[2118] ), .B1(_04620_ ), .B2(_02339_ ), .ZN(_04625_ ) );
AOI21_X1 _19134_ ( .A(fanout_net_59 ), .B1(_04624_ ), .B2(_04625_ ), .ZN(_01706_ ) );
BUF_X4 _19135_ ( .A(_09953_ ), .Z(_04626_ ) );
NAND4_X1 _19136_ ( .A1(_04626_ ), .A2(_09961_ ), .A3(_09979_ ), .A4(_03978_ ), .ZN(_04627_ ) );
OAI21_X1 _19137_ ( .A(\u_lsu.pmem[2117] ), .B1(_04620_ ), .B2(_02339_ ), .ZN(_04628_ ) );
AOI21_X1 _19138_ ( .A(fanout_net_59 ), .B1(_04627_ ), .B2(_04628_ ), .ZN(_01707_ ) );
NAND4_X1 _19139_ ( .A1(_04626_ ), .A2(_09966_ ), .A3(_09979_ ), .A4(_03978_ ), .ZN(_04629_ ) );
OAI21_X1 _19140_ ( .A(\u_lsu.pmem[2116] ), .B1(_04620_ ), .B2(_02337_ ), .ZN(_04630_ ) );
AOI21_X1 _19141_ ( .A(fanout_net_59 ), .B1(_04629_ ), .B2(_04630_ ), .ZN(_01708_ ) );
NAND4_X1 _19142_ ( .A1(_04626_ ), .A2(_09970_ ), .A3(_09979_ ), .A4(_09879_ ), .ZN(_04631_ ) );
OAI21_X1 _19143_ ( .A(\u_lsu.pmem[2115] ), .B1(_04620_ ), .B2(_02337_ ), .ZN(_04632_ ) );
AOI21_X1 _19144_ ( .A(fanout_net_59 ), .B1(_04631_ ), .B2(_04632_ ), .ZN(_01709_ ) );
OAI21_X1 _19145_ ( .A(\u_lsu.pmem[4163] ), .B1(_04583_ ), .B2(_09949_ ), .ZN(_04633_ ) );
NAND4_X1 _19146_ ( .A1(_09970_ ), .A2(_04585_ ), .A3(_04556_ ), .A4(_11159_ ), .ZN(_04634_ ) );
AOI21_X1 _19147_ ( .A(fanout_net_59 ), .B1(_04633_ ), .B2(_04634_ ), .ZN(_01710_ ) );
NAND4_X1 _19148_ ( .A1(_04626_ ), .A2(_09974_ ), .A3(_09979_ ), .A4(_09879_ ), .ZN(_04635_ ) );
OAI21_X1 _19149_ ( .A(\u_lsu.pmem[2114] ), .B1(_04620_ ), .B2(_02337_ ), .ZN(_04636_ ) );
AOI21_X1 _19150_ ( .A(fanout_net_59 ), .B1(_04635_ ), .B2(_04636_ ), .ZN(_01711_ ) );
NAND4_X1 _19151_ ( .A1(_04626_ ), .A2(_09978_ ), .A3(_09540_ ), .A4(_09879_ ), .ZN(_04637_ ) );
OAI21_X1 _19152_ ( .A(\u_lsu.pmem[2113] ), .B1(_04620_ ), .B2(_02337_ ), .ZN(_04638_ ) );
AOI21_X1 _19153_ ( .A(fanout_net_59 ), .B1(_04637_ ), .B2(_04638_ ), .ZN(_01712_ ) );
NAND4_X1 _19154_ ( .A1(_04626_ ), .A2(_09982_ ), .A3(_09540_ ), .A4(_09879_ ), .ZN(_04639_ ) );
OAI21_X1 _19155_ ( .A(\u_lsu.pmem[2112] ), .B1(_04620_ ), .B2(_02337_ ), .ZN(_04640_ ) );
AOI21_X1 _19156_ ( .A(fanout_net_59 ), .B1(_04639_ ), .B2(_04640_ ), .ZN(_01713_ ) );
NAND4_X1 _19157_ ( .A1(_09987_ ), .A2(_04574_ ), .A3(_04560_ ), .A4(_04567_ ), .ZN(_04641_ ) );
OAI21_X1 _19158_ ( .A(\u_lsu.pmem[2087] ), .B1(_04620_ ), .B2(_02363_ ), .ZN(_04642_ ) );
AOI21_X1 _19159_ ( .A(fanout_net_59 ), .B1(_04641_ ), .B2(_04642_ ), .ZN(_01714_ ) );
NAND4_X1 _19160_ ( .A1(_09994_ ), .A2(_04574_ ), .A3(_04560_ ), .A4(_04567_ ), .ZN(_04643_ ) );
OAI21_X1 _19161_ ( .A(\u_lsu.pmem[2086] ), .B1(_04620_ ), .B2(_02363_ ), .ZN(_04644_ ) );
AOI21_X1 _19162_ ( .A(fanout_net_59 ), .B1(_04643_ ), .B2(_04644_ ), .ZN(_01715_ ) );
NAND4_X1 _19163_ ( .A1(_09997_ ), .A2(_04574_ ), .A3(_04560_ ), .A4(_04567_ ), .ZN(_04645_ ) );
BUF_X4 _19164_ ( .A(_04571_ ), .Z(_04646_ ) );
OAI21_X1 _19165_ ( .A(\u_lsu.pmem[2085] ), .B1(_04646_ ), .B2(_02363_ ), .ZN(_04647_ ) );
AOI21_X1 _19166_ ( .A(fanout_net_59 ), .B1(_04645_ ), .B2(_04647_ ), .ZN(_01716_ ) );
NOR2_X1 _19167_ ( .A1(_09141_ ), .A2(_02362_ ), .ZN(_04648_ ) );
OAI21_X1 _19168_ ( .A(_09109_ ), .B1(_04648_ ), .B2(\u_lsu.pmem[2084] ), .ZN(_04649_ ) );
AOI21_X1 _19169_ ( .A(_04649_ ), .B1(_09149_ ), .B2(_04648_ ), .ZN(_01717_ ) );
NAND2_X1 _19170_ ( .A1(_04648_ ), .A2(_03114_ ), .ZN(_04650_ ) );
OAI21_X1 _19171_ ( .A(\u_lsu.pmem[2083] ), .B1(_04646_ ), .B2(_02362_ ), .ZN(_04651_ ) );
AOI21_X1 _19172_ ( .A(fanout_net_59 ), .B1(_04650_ ), .B2(_04651_ ), .ZN(_01718_ ) );
NAND2_X1 _19173_ ( .A1(_04648_ ), .A2(_03145_ ), .ZN(_04652_ ) );
OAI21_X1 _19174_ ( .A(\u_lsu.pmem[2082] ), .B1(_04646_ ), .B2(_02362_ ), .ZN(_04653_ ) );
AOI21_X1 _19175_ ( .A(fanout_net_59 ), .B1(_04652_ ), .B2(_04653_ ), .ZN(_01719_ ) );
NAND2_X1 _19176_ ( .A1(_04648_ ), .A2(_03174_ ), .ZN(_04654_ ) );
OAI21_X1 _19177_ ( .A(\u_lsu.pmem[2081] ), .B1(_04646_ ), .B2(_02362_ ), .ZN(_04655_ ) );
AOI21_X1 _19178_ ( .A(fanout_net_59 ), .B1(_04654_ ), .B2(_04655_ ), .ZN(_01720_ ) );
OAI21_X1 _19179_ ( .A(\u_lsu.pmem[4162] ), .B1(_04583_ ), .B2(_09949_ ), .ZN(_04656_ ) );
NAND4_X1 _19180_ ( .A1(_09974_ ), .A2(_04585_ ), .A3(_04556_ ), .A4(_11159_ ), .ZN(_04657_ ) );
AOI21_X1 _19181_ ( .A(fanout_net_59 ), .B1(_04656_ ), .B2(_04657_ ), .ZN(_01721_ ) );
BUF_X4 _19182_ ( .A(_10578_ ), .Z(_04658_ ) );
NAND4_X1 _19183_ ( .A1(_10021_ ), .A2(_04574_ ), .A3(_04658_ ), .A4(_04567_ ), .ZN(_04659_ ) );
OAI21_X1 _19184_ ( .A(\u_lsu.pmem[2080] ), .B1(_04646_ ), .B2(_02362_ ), .ZN(_04660_ ) );
AOI21_X1 _19185_ ( .A(fanout_net_59 ), .B1(_04659_ ), .B2(_04660_ ), .ZN(_01722_ ) );
NAND4_X1 _19186_ ( .A1(_02387_ ), .A2(_11423_ ), .A3(_10071_ ), .A4(_09607_ ), .ZN(_04661_ ) );
OAI21_X1 _19187_ ( .A(\u_lsu.pmem[2055] ), .B1(_02390_ ), .B2(_04013_ ), .ZN(_04662_ ) );
AOI21_X1 _19188_ ( .A(fanout_net_59 ), .B1(_04661_ ), .B2(_04662_ ), .ZN(_01723_ ) );
NAND4_X1 _19189_ ( .A1(_02387_ ), .A2(_09658_ ), .A3(_10071_ ), .A4(_09607_ ), .ZN(_04663_ ) );
OAI21_X1 _19190_ ( .A(\u_lsu.pmem[2054] ), .B1(_02390_ ), .B2(_04013_ ), .ZN(_04664_ ) );
AOI21_X1 _19191_ ( .A(fanout_net_59 ), .B1(_04663_ ), .B2(_04664_ ), .ZN(_01724_ ) );
NAND4_X1 _19192_ ( .A1(_02387_ ), .A2(_09713_ ), .A3(_10071_ ), .A4(_09607_ ), .ZN(_04665_ ) );
OAI21_X1 _19193_ ( .A(\u_lsu.pmem[2053] ), .B1(_02390_ ), .B2(_04013_ ), .ZN(_04666_ ) );
AOI21_X1 _19194_ ( .A(fanout_net_59 ), .B1(_04665_ ), .B2(_04666_ ), .ZN(_01725_ ) );
NAND4_X1 _19195_ ( .A1(_02387_ ), .A2(_09514_ ), .A3(_10071_ ), .A4(_09607_ ), .ZN(_04667_ ) );
OAI21_X1 _19196_ ( .A(\u_lsu.pmem[2052] ), .B1(_02389_ ), .B2(_04013_ ), .ZN(_04668_ ) );
AOI21_X1 _19197_ ( .A(fanout_net_59 ), .B1(_04667_ ), .B2(_04668_ ), .ZN(_01726_ ) );
BUF_X4 _19198_ ( .A(_09133_ ), .Z(_04669_ ) );
NAND4_X1 _19199_ ( .A1(_04669_ ), .A2(_10456_ ), .A3(_10071_ ), .A4(_09607_ ), .ZN(_04670_ ) );
BUF_X4 _19200_ ( .A(_10041_ ), .Z(_04671_ ) );
OAI21_X1 _19201_ ( .A(\u_lsu.pmem[2051] ), .B1(_02389_ ), .B2(_04671_ ), .ZN(_04672_ ) );
AOI21_X1 _19202_ ( .A(fanout_net_59 ), .B1(_04670_ ), .B2(_04672_ ), .ZN(_01727_ ) );
NAND4_X1 _19203_ ( .A1(_11021_ ), .A2(_03909_ ), .A3(_04454_ ), .A4(_04567_ ), .ZN(_04673_ ) );
OAI21_X1 _19204_ ( .A(\u_lsu.pmem[2050] ), .B1(_02389_ ), .B2(_04671_ ), .ZN(_04674_ ) );
AOI21_X1 _19205_ ( .A(fanout_net_59 ), .B1(_04673_ ), .B2(_04674_ ), .ZN(_01728_ ) );
NAND4_X1 _19206_ ( .A1(_04669_ ), .A2(_09544_ ), .A3(_10071_ ), .A4(_09607_ ), .ZN(_04675_ ) );
OAI21_X1 _19207_ ( .A(\u_lsu.pmem[2049] ), .B1(_02389_ ), .B2(_04671_ ), .ZN(_04676_ ) );
AOI21_X1 _19208_ ( .A(fanout_net_59 ), .B1(_04675_ ), .B2(_04676_ ), .ZN(_01729_ ) );
NAND4_X1 _19209_ ( .A1(_04669_ ), .A2(_10467_ ), .A3(_10071_ ), .A4(_09607_ ), .ZN(_04677_ ) );
OAI21_X1 _19210_ ( .A(\u_lsu.pmem[2048] ), .B1(_02389_ ), .B2(_04671_ ), .ZN(_04678_ ) );
AOI21_X1 _19211_ ( .A(fanout_net_60 ), .B1(_04677_ ), .B2(_04678_ ), .ZN(_01730_ ) );
NOR2_X1 _19212_ ( .A1(_10033_ ), .A2(_02410_ ), .ZN(_04679_ ) );
NOR2_X1 _19213_ ( .A1(_04679_ ), .A2(\u_lsu.pmem[2023] ), .ZN(_04680_ ) );
AOI211_X1 _19214_ ( .A(fanout_net_60 ), .B(_04680_ ), .C1(_04216_ ), .C2(_04679_ ), .ZN(_01731_ ) );
OAI21_X1 _19215_ ( .A(\u_lsu.pmem[4161] ), .B1(_04583_ ), .B2(_09949_ ), .ZN(_04681_ ) );
NAND4_X1 _19216_ ( .A1(_09978_ ), .A2(_04585_ ), .A3(_04556_ ), .A4(_11159_ ), .ZN(_04682_ ) );
AOI21_X1 _19217_ ( .A(fanout_net_60 ), .B1(_04681_ ), .B2(_04682_ ), .ZN(_01732_ ) );
NAND4_X1 _19218_ ( .A1(_10062_ ), .A2(_03909_ ), .A3(_04454_ ), .A4(_04567_ ), .ZN(_04683_ ) );
OAI21_X1 _19219_ ( .A(\u_lsu.pmem[2022] ), .B1(_04646_ ), .B2(_02411_ ), .ZN(_04684_ ) );
AOI21_X1 _19220_ ( .A(fanout_net_60 ), .B1(_04683_ ), .B2(_04684_ ), .ZN(_01733_ ) );
BUF_X8 _19221_ ( .A(_09442_ ), .Z(_04685_ ) );
BUF_X4 _19222_ ( .A(_04685_ ), .Z(_04686_ ) );
NAND4_X1 _19223_ ( .A1(_10075_ ), .A2(_03909_ ), .A3(_04454_ ), .A4(_04686_ ), .ZN(_04687_ ) );
OAI21_X1 _19224_ ( .A(\u_lsu.pmem[2021] ), .B1(_04646_ ), .B2(_02411_ ), .ZN(_04688_ ) );
AOI21_X1 _19225_ ( .A(fanout_net_60 ), .B1(_04687_ ), .B2(_04688_ ), .ZN(_01734_ ) );
BUF_X4 _19226_ ( .A(_03020_ ), .Z(_04689_ ) );
NAND4_X1 _19227_ ( .A1(_10079_ ), .A2(_04689_ ), .A3(_04454_ ), .A4(_04686_ ), .ZN(_04690_ ) );
OAI21_X1 _19228_ ( .A(\u_lsu.pmem[2020] ), .B1(_04646_ ), .B2(_02410_ ), .ZN(_04691_ ) );
AOI21_X1 _19229_ ( .A(fanout_net_60 ), .B1(_04690_ ), .B2(_04691_ ), .ZN(_01735_ ) );
NAND4_X1 _19230_ ( .A1(_10084_ ), .A2(_04689_ ), .A3(_04454_ ), .A4(_04686_ ), .ZN(_04692_ ) );
OAI21_X1 _19231_ ( .A(\u_lsu.pmem[2019] ), .B1(_04646_ ), .B2(_02410_ ), .ZN(_04693_ ) );
AOI21_X1 _19232_ ( .A(fanout_net_60 ), .B1(_04692_ ), .B2(_04693_ ), .ZN(_01736_ ) );
NAND4_X1 _19233_ ( .A1(_10088_ ), .A2(_04689_ ), .A3(_04454_ ), .A4(_04686_ ), .ZN(_04694_ ) );
OAI21_X1 _19234_ ( .A(\u_lsu.pmem[2018] ), .B1(_04646_ ), .B2(_02410_ ), .ZN(_04695_ ) );
AOI21_X1 _19235_ ( .A(fanout_net_60 ), .B1(_04694_ ), .B2(_04695_ ), .ZN(_01737_ ) );
NAND4_X1 _19236_ ( .A1(_10094_ ), .A2(_04689_ ), .A3(_04454_ ), .A4(_04686_ ), .ZN(_04696_ ) );
BUF_X4 _19237_ ( .A(_04571_ ), .Z(_04697_ ) );
OAI21_X1 _19238_ ( .A(\u_lsu.pmem[2017] ), .B1(_04697_ ), .B2(_02410_ ), .ZN(_04698_ ) );
AOI21_X1 _19239_ ( .A(fanout_net_60 ), .B1(_04696_ ), .B2(_04698_ ), .ZN(_01738_ ) );
NAND4_X1 _19240_ ( .A1(_10098_ ), .A2(_04689_ ), .A3(_04454_ ), .A4(_04686_ ), .ZN(_04699_ ) );
OAI21_X1 _19241_ ( .A(\u_lsu.pmem[2016] ), .B1(_04697_ ), .B2(_02410_ ), .ZN(_04700_ ) );
AOI21_X1 _19242_ ( .A(fanout_net_60 ), .B1(_04699_ ), .B2(_04700_ ), .ZN(_01739_ ) );
NAND4_X1 _19243_ ( .A1(_04626_ ), .A2(_02486_ ), .A3(_09914_ ), .A4(_10104_ ), .ZN(_04701_ ) );
OAI21_X1 _19244_ ( .A(\u_lsu.pmem[1991] ), .B1(_04697_ ), .B2(_02435_ ), .ZN(_04702_ ) );
AOI21_X1 _19245_ ( .A(fanout_net_60 ), .B1(_04701_ ), .B2(_04702_ ), .ZN(_01740_ ) );
NAND4_X1 _19246_ ( .A1(_10117_ ), .A2(_04689_ ), .A3(_04454_ ), .A4(_04686_ ), .ZN(_04703_ ) );
OAI21_X1 _19247_ ( .A(\u_lsu.pmem[1990] ), .B1(_04697_ ), .B2(_02435_ ), .ZN(_04704_ ) );
AOI21_X1 _19248_ ( .A(fanout_net_60 ), .B1(_04703_ ), .B2(_04704_ ), .ZN(_01741_ ) );
BUF_X4 _19249_ ( .A(_03326_ ), .Z(_04705_ ) );
NAND4_X1 _19250_ ( .A1(_10121_ ), .A2(_04689_ ), .A3(_04705_ ), .A4(_04686_ ), .ZN(_04706_ ) );
OAI21_X1 _19251_ ( .A(\u_lsu.pmem[1989] ), .B1(_04697_ ), .B2(_02434_ ), .ZN(_04707_ ) );
AOI21_X1 _19252_ ( .A(fanout_net_60 ), .B1(_04706_ ), .B2(_04707_ ), .ZN(_01742_ ) );
NAND4_X1 _19253_ ( .A1(_09715_ ), .A2(_04574_ ), .A3(_04705_ ), .A4(_04097_ ), .ZN(_04708_ ) );
OAI21_X1 _19254_ ( .A(\u_lsu.pmem[4358] ), .B1(_04071_ ), .B2(_09468_ ), .ZN(_04709_ ) );
AOI21_X1 _19255_ ( .A(fanout_net_60 ), .B1(_04708_ ), .B2(_04709_ ), .ZN(_01743_ ) );
OAI21_X1 _19256_ ( .A(\u_lsu.pmem[4160] ), .B1(_04583_ ), .B2(_09949_ ), .ZN(_04710_ ) );
NAND4_X1 _19257_ ( .A1(_09982_ ), .A2(_04585_ ), .A3(_04556_ ), .A4(_11159_ ), .ZN(_04711_ ) );
AOI21_X1 _19258_ ( .A(fanout_net_60 ), .B1(_04710_ ), .B2(_04711_ ), .ZN(_01744_ ) );
NAND4_X1 _19259_ ( .A1(_10125_ ), .A2(_04689_ ), .A3(_04705_ ), .A4(_04686_ ), .ZN(_04712_ ) );
OAI21_X1 _19260_ ( .A(\u_lsu.pmem[1988] ), .B1(_04697_ ), .B2(_02434_ ), .ZN(_04713_ ) );
AOI21_X1 _19261_ ( .A(fanout_net_60 ), .B1(_04712_ ), .B2(_04713_ ), .ZN(_01745_ ) );
NAND4_X1 _19262_ ( .A1(_10131_ ), .A2(_04689_ ), .A3(_04705_ ), .A4(_04686_ ), .ZN(_04714_ ) );
OAI21_X1 _19263_ ( .A(\u_lsu.pmem[1987] ), .B1(_04697_ ), .B2(_02434_ ), .ZN(_04715_ ) );
AOI21_X1 _19264_ ( .A(fanout_net_60 ), .B1(_04714_ ), .B2(_04715_ ), .ZN(_01746_ ) );
BUF_X4 _19265_ ( .A(_04685_ ), .Z(_04716_ ) );
NAND4_X1 _19266_ ( .A1(_10135_ ), .A2(_04689_ ), .A3(_04705_ ), .A4(_04716_ ), .ZN(_04717_ ) );
OAI21_X1 _19267_ ( .A(\u_lsu.pmem[1986] ), .B1(_04697_ ), .B2(_02434_ ), .ZN(_04718_ ) );
AOI21_X1 _19268_ ( .A(fanout_net_60 ), .B1(_04717_ ), .B2(_04718_ ), .ZN(_01747_ ) );
BUF_X4 _19269_ ( .A(_03020_ ), .Z(_04719_ ) );
NAND4_X1 _19270_ ( .A1(_10138_ ), .A2(_04719_ ), .A3(_04705_ ), .A4(_04716_ ), .ZN(_04720_ ) );
OAI21_X1 _19271_ ( .A(\u_lsu.pmem[1985] ), .B1(_04697_ ), .B2(_02434_ ), .ZN(_04721_ ) );
AOI21_X1 _19272_ ( .A(fanout_net_60 ), .B1(_04720_ ), .B2(_04721_ ), .ZN(_01748_ ) );
NAND4_X1 _19273_ ( .A1(_10144_ ), .A2(_04719_ ), .A3(_04705_ ), .A4(_04716_ ), .ZN(_04722_ ) );
OAI21_X1 _19274_ ( .A(\u_lsu.pmem[1984] ), .B1(_04697_ ), .B2(_02434_ ), .ZN(_04723_ ) );
AOI21_X1 _19275_ ( .A(fanout_net_60 ), .B1(_04722_ ), .B2(_04723_ ), .ZN(_01749_ ) );
NAND4_X1 _19276_ ( .A1(_10148_ ), .A2(_04719_ ), .A3(_04705_ ), .A4(_04716_ ), .ZN(_04724_ ) );
BUF_X4 _19277_ ( .A(_04571_ ), .Z(_04725_ ) );
OAI21_X1 _19278_ ( .A(\u_lsu.pmem[1959] ), .B1(_04725_ ), .B2(_02460_ ), .ZN(_04726_ ) );
AOI21_X1 _19279_ ( .A(fanout_net_60 ), .B1(_04724_ ), .B2(_04726_ ), .ZN(_01750_ ) );
NAND4_X1 _19280_ ( .A1(_10156_ ), .A2(_04719_ ), .A3(_04705_ ), .A4(_04716_ ), .ZN(_04727_ ) );
OAI21_X1 _19281_ ( .A(\u_lsu.pmem[1958] ), .B1(_04725_ ), .B2(_02460_ ), .ZN(_04728_ ) );
AOI21_X1 _19282_ ( .A(fanout_net_60 ), .B1(_04727_ ), .B2(_04728_ ), .ZN(_01751_ ) );
NAND4_X1 _19283_ ( .A1(_10160_ ), .A2(_04719_ ), .A3(_04705_ ), .A4(_04716_ ), .ZN(_04729_ ) );
OAI21_X1 _19284_ ( .A(\u_lsu.pmem[1957] ), .B1(_04725_ ), .B2(_02459_ ), .ZN(_04730_ ) );
AOI21_X1 _19285_ ( .A(fanout_net_60 ), .B1(_04729_ ), .B2(_04730_ ), .ZN(_01752_ ) );
BUF_X8 _19286_ ( .A(_09455_ ), .Z(_04731_ ) );
BUF_X4 _19287_ ( .A(_04731_ ), .Z(_04732_ ) );
NAND4_X1 _19288_ ( .A1(_10166_ ), .A2(_04719_ ), .A3(_04732_ ), .A4(_04716_ ), .ZN(_04733_ ) );
OAI21_X1 _19289_ ( .A(\u_lsu.pmem[1956] ), .B1(_04725_ ), .B2(_02459_ ), .ZN(_04734_ ) );
AOI21_X1 _19290_ ( .A(fanout_net_60 ), .B1(_04733_ ), .B2(_04734_ ), .ZN(_01753_ ) );
NAND4_X1 _19291_ ( .A1(_10169_ ), .A2(_04719_ ), .A3(_04732_ ), .A4(_04716_ ), .ZN(_04735_ ) );
OAI21_X1 _19292_ ( .A(\u_lsu.pmem[1955] ), .B1(_04725_ ), .B2(_02459_ ), .ZN(_04736_ ) );
AOI21_X1 _19293_ ( .A(fanout_net_60 ), .B1(_04735_ ), .B2(_04736_ ), .ZN(_01754_ ) );
NAND4_X1 _19294_ ( .A1(_09987_ ), .A2(_04574_ ), .A3(_04732_ ), .A4(_04097_ ), .ZN(_04737_ ) );
OAI21_X1 _19295_ ( .A(\u_lsu.pmem[4135] ), .B1(_04071_ ), .B2(_09991_ ), .ZN(_04738_ ) );
AOI21_X1 _19296_ ( .A(fanout_net_60 ), .B1(_04737_ ), .B2(_04738_ ), .ZN(_01755_ ) );
NAND4_X1 _19297_ ( .A1(_10172_ ), .A2(_04719_ ), .A3(_04732_ ), .A4(_04716_ ), .ZN(_04739_ ) );
OAI21_X1 _19298_ ( .A(\u_lsu.pmem[1954] ), .B1(_04725_ ), .B2(_02459_ ), .ZN(_04740_ ) );
AOI21_X1 _19299_ ( .A(fanout_net_60 ), .B1(_04739_ ), .B2(_04740_ ), .ZN(_01756_ ) );
NAND4_X1 _19300_ ( .A1(_10176_ ), .A2(_04719_ ), .A3(_04732_ ), .A4(_04716_ ), .ZN(_04741_ ) );
OAI21_X1 _19301_ ( .A(\u_lsu.pmem[1953] ), .B1(_04725_ ), .B2(_02459_ ), .ZN(_04742_ ) );
AOI21_X1 _19302_ ( .A(fanout_net_60 ), .B1(_04741_ ), .B2(_04742_ ), .ZN(_01757_ ) );
NAND3_X1 _19303_ ( .A1(_04009_ ), .A2(_03203_ ), .A3(_02458_ ), .ZN(_04743_ ) );
OAI21_X1 _19304_ ( .A(\u_lsu.pmem[1952] ), .B1(_04725_ ), .B2(_02459_ ), .ZN(_04744_ ) );
AOI21_X1 _19305_ ( .A(fanout_net_60 ), .B1(_04743_ ), .B2(_04744_ ), .ZN(_01758_ ) );
BUF_X4 _19306_ ( .A(_04685_ ), .Z(_04745_ ) );
NAND4_X1 _19307_ ( .A1(_02483_ ), .A2(_09603_ ), .A3(_02500_ ), .A4(_04745_ ), .ZN(_04746_ ) );
OAI21_X1 _19308_ ( .A(\u_lsu.pmem[1927] ), .B1(_02489_ ), .B2(_04410_ ), .ZN(_04747_ ) );
AOI21_X1 _19309_ ( .A(fanout_net_60 ), .B1(_04746_ ), .B2(_04747_ ), .ZN(_01759_ ) );
NAND4_X1 _19310_ ( .A1(_02483_ ), .A2(_09658_ ), .A3(_02500_ ), .A4(_04745_ ), .ZN(_04748_ ) );
OAI21_X1 _19311_ ( .A(\u_lsu.pmem[1926] ), .B1(_02488_ ), .B2(_04410_ ), .ZN(_04749_ ) );
AOI21_X1 _19312_ ( .A(fanout_net_61 ), .B1(_04748_ ), .B2(_04749_ ), .ZN(_01760_ ) );
NAND4_X1 _19313_ ( .A1(_02483_ ), .A2(_09713_ ), .A3(_03436_ ), .A4(_04745_ ), .ZN(_04750_ ) );
OAI21_X1 _19314_ ( .A(\u_lsu.pmem[1925] ), .B1(_02488_ ), .B2(_04410_ ), .ZN(_04751_ ) );
AOI21_X1 _19315_ ( .A(fanout_net_61 ), .B1(_04750_ ), .B2(_04751_ ), .ZN(_01761_ ) );
NAND4_X1 _19316_ ( .A1(_09602_ ), .A2(_09514_ ), .A3(_03436_ ), .A4(_04745_ ), .ZN(_04752_ ) );
BUF_X4 _19317_ ( .A(_04265_ ), .Z(_04753_ ) );
OAI21_X1 _19318_ ( .A(\u_lsu.pmem[1924] ), .B1(_02488_ ), .B2(_04753_ ), .ZN(_04754_ ) );
AOI21_X1 _19319_ ( .A(fanout_net_61 ), .B1(_04752_ ), .B2(_04754_ ), .ZN(_01762_ ) );
NAND4_X1 _19320_ ( .A1(_09602_ ), .A2(_10456_ ), .A3(_03436_ ), .A4(_04745_ ), .ZN(_04755_ ) );
OAI21_X1 _19321_ ( .A(\u_lsu.pmem[1923] ), .B1(_02488_ ), .B2(_04753_ ), .ZN(_04756_ ) );
AOI21_X1 _19322_ ( .A(fanout_net_61 ), .B1(_04755_ ), .B2(_04756_ ), .ZN(_01763_ ) );
OAI21_X1 _19323_ ( .A(\u_lsu.pmem[1922] ), .B1(_02489_ ), .B2(_04593_ ), .ZN(_04757_ ) );
NAND4_X1 _19324_ ( .A1(_09874_ ), .A2(_03107_ ), .A3(_04556_ ), .A4(_04595_ ), .ZN(_04758_ ) );
AOI21_X1 _19325_ ( .A(fanout_net_61 ), .B1(_04757_ ), .B2(_04758_ ), .ZN(_01764_ ) );
NAND4_X1 _19326_ ( .A1(_09602_ ), .A2(_09544_ ), .A3(_03436_ ), .A4(_04745_ ), .ZN(_04759_ ) );
OAI21_X1 _19327_ ( .A(\u_lsu.pmem[1921] ), .B1(_02488_ ), .B2(_04753_ ), .ZN(_04760_ ) );
AOI21_X1 _19328_ ( .A(fanout_net_61 ), .B1(_04759_ ), .B2(_04760_ ), .ZN(_01765_ ) );
NAND4_X1 _19329_ ( .A1(_09994_ ), .A2(_04574_ ), .A3(_04732_ ), .A4(_04097_ ), .ZN(_04761_ ) );
OAI21_X1 _19330_ ( .A(\u_lsu.pmem[4134] ), .B1(_04071_ ), .B2(_09991_ ), .ZN(_04762_ ) );
AOI21_X1 _19331_ ( .A(fanout_net_61 ), .B1(_04761_ ), .B2(_04762_ ), .ZN(_01766_ ) );
NAND4_X1 _19332_ ( .A1(_09602_ ), .A2(_10467_ ), .A3(_03436_ ), .A4(_04745_ ), .ZN(_04763_ ) );
OAI21_X1 _19333_ ( .A(\u_lsu.pmem[1920] ), .B1(_02488_ ), .B2(_04753_ ), .ZN(_04764_ ) );
AOI21_X1 _19334_ ( .A(fanout_net_61 ), .B1(_04763_ ), .B2(_04764_ ), .ZN(_01767_ ) );
NAND3_X1 _19335_ ( .A1(_04009_ ), .A2(_11138_ ), .A3(_02509_ ), .ZN(_04765_ ) );
OAI21_X1 _19336_ ( .A(\u_lsu.pmem[1895] ), .B1(_04725_ ), .B2(_02512_ ), .ZN(_04766_ ) );
AOI21_X1 _19337_ ( .A(fanout_net_61 ), .B1(_04765_ ), .B2(_04766_ ), .ZN(_01768_ ) );
NAND3_X1 _19338_ ( .A1(_04009_ ), .A2(_11145_ ), .A3(_02509_ ), .ZN(_04767_ ) );
OAI21_X1 _19339_ ( .A(\u_lsu.pmem[1894] ), .B1(_04725_ ), .B2(_02512_ ), .ZN(_04768_ ) );
AOI21_X1 _19340_ ( .A(fanout_net_61 ), .B1(_04767_ ), .B2(_04768_ ), .ZN(_01769_ ) );
NAND3_X1 _19341_ ( .A1(_04009_ ), .A2(_11148_ ), .A3(_02509_ ), .ZN(_04769_ ) );
BUF_X4 _19342_ ( .A(_04571_ ), .Z(_04770_ ) );
OAI21_X1 _19343_ ( .A(\u_lsu.pmem[1893] ), .B1(_04770_ ), .B2(_02511_ ), .ZN(_04771_ ) );
AOI21_X1 _19344_ ( .A(fanout_net_61 ), .B1(_04769_ ), .B2(_04771_ ), .ZN(_01770_ ) );
BUF_X4 _19345_ ( .A(_04008_ ), .Z(_04772_ ) );
NAND3_X1 _19346_ ( .A1(_04772_ ), .A2(_03084_ ), .A3(_02509_ ), .ZN(_04773_ ) );
OAI21_X1 _19347_ ( .A(\u_lsu.pmem[1892] ), .B1(_04770_ ), .B2(_02511_ ), .ZN(_04774_ ) );
AOI21_X1 _19348_ ( .A(fanout_net_61 ), .B1(_04773_ ), .B2(_04774_ ), .ZN(_01771_ ) );
NAND3_X1 _19349_ ( .A1(_04772_ ), .A2(_03114_ ), .A3(_02509_ ), .ZN(_04775_ ) );
OAI21_X1 _19350_ ( .A(\u_lsu.pmem[1891] ), .B1(_04770_ ), .B2(_02511_ ), .ZN(_04776_ ) );
AOI21_X1 _19351_ ( .A(fanout_net_61 ), .B1(_04775_ ), .B2(_04776_ ), .ZN(_01772_ ) );
NAND3_X1 _19352_ ( .A1(_04772_ ), .A2(_03145_ ), .A3(_02509_ ), .ZN(_04777_ ) );
OAI21_X1 _19353_ ( .A(\u_lsu.pmem[1890] ), .B1(_04770_ ), .B2(_02511_ ), .ZN(_04778_ ) );
AOI21_X1 _19354_ ( .A(fanout_net_61 ), .B1(_04777_ ), .B2(_04778_ ), .ZN(_01773_ ) );
NAND3_X1 _19355_ ( .A1(_04772_ ), .A2(_03174_ ), .A3(_02509_ ), .ZN(_04779_ ) );
OAI21_X1 _19356_ ( .A(\u_lsu.pmem[1889] ), .B1(_04770_ ), .B2(_02511_ ), .ZN(_04780_ ) );
AOI21_X1 _19357_ ( .A(fanout_net_61 ), .B1(_04779_ ), .B2(_04780_ ), .ZN(_01774_ ) );
NAND3_X1 _19358_ ( .A1(_04772_ ), .A2(_03203_ ), .A3(_02509_ ), .ZN(_04781_ ) );
OAI21_X1 _19359_ ( .A(\u_lsu.pmem[1888] ), .B1(_04770_ ), .B2(_02511_ ), .ZN(_04782_ ) );
AOI21_X1 _19360_ ( .A(fanout_net_61 ), .B1(_04781_ ), .B2(_04782_ ), .ZN(_01775_ ) );
NAND3_X1 _19361_ ( .A1(_04772_ ), .A2(_11138_ ), .A3(_02535_ ), .ZN(_04783_ ) );
OAI21_X1 _19362_ ( .A(\u_lsu.pmem[1863] ), .B1(_04770_ ), .B2(_02538_ ), .ZN(_04784_ ) );
AOI21_X1 _19363_ ( .A(fanout_net_61 ), .B1(_04783_ ), .B2(_04784_ ), .ZN(_01776_ ) );
NAND4_X1 _19364_ ( .A1(_09997_ ), .A2(_04574_ ), .A3(_04732_ ), .A4(_04097_ ), .ZN(_04785_ ) );
OAI21_X1 _19365_ ( .A(\u_lsu.pmem[4133] ), .B1(_04071_ ), .B2(_09991_ ), .ZN(_04786_ ) );
AOI21_X1 _19366_ ( .A(fanout_net_61 ), .B1(_04785_ ), .B2(_04786_ ), .ZN(_01777_ ) );
NAND3_X1 _19367_ ( .A1(_04772_ ), .A2(_11145_ ), .A3(_02535_ ), .ZN(_04787_ ) );
OAI21_X1 _19368_ ( .A(\u_lsu.pmem[1862] ), .B1(_04770_ ), .B2(_02538_ ), .ZN(_04788_ ) );
AOI21_X1 _19369_ ( .A(fanout_net_61 ), .B1(_04787_ ), .B2(_04788_ ), .ZN(_01778_ ) );
NAND3_X1 _19370_ ( .A1(_04772_ ), .A2(_11148_ ), .A3(_02535_ ), .ZN(_04789_ ) );
OAI21_X1 _19371_ ( .A(\u_lsu.pmem[1861] ), .B1(_04770_ ), .B2(_02537_ ), .ZN(_04790_ ) );
AOI21_X1 _19372_ ( .A(fanout_net_61 ), .B1(_04789_ ), .B2(_04790_ ), .ZN(_01779_ ) );
NAND3_X1 _19373_ ( .A1(_04772_ ), .A2(_03084_ ), .A3(_02535_ ), .ZN(_04791_ ) );
OAI21_X1 _19374_ ( .A(\u_lsu.pmem[1860] ), .B1(_04770_ ), .B2(_02537_ ), .ZN(_04792_ ) );
AOI21_X1 _19375_ ( .A(fanout_net_61 ), .B1(_04791_ ), .B2(_04792_ ), .ZN(_01780_ ) );
NAND3_X1 _19376_ ( .A1(_04772_ ), .A2(_03114_ ), .A3(_02535_ ), .ZN(_04793_ ) );
BUF_X4 _19377_ ( .A(_04571_ ), .Z(_04794_ ) );
OAI21_X1 _19378_ ( .A(\u_lsu.pmem[1859] ), .B1(_04794_ ), .B2(_02537_ ), .ZN(_04795_ ) );
AOI21_X1 _19379_ ( .A(fanout_net_61 ), .B1(_04793_ ), .B2(_04795_ ), .ZN(_01781_ ) );
BUF_X4 _19380_ ( .A(_04008_ ), .Z(_04796_ ) );
NAND3_X1 _19381_ ( .A1(_04796_ ), .A2(_03145_ ), .A3(_02535_ ), .ZN(_04797_ ) );
OAI21_X1 _19382_ ( .A(\u_lsu.pmem[1858] ), .B1(_04794_ ), .B2(_02537_ ), .ZN(_04798_ ) );
AOI21_X1 _19383_ ( .A(fanout_net_61 ), .B1(_04797_ ), .B2(_04798_ ), .ZN(_01782_ ) );
NAND3_X1 _19384_ ( .A1(_04796_ ), .A2(_03174_ ), .A3(_02535_ ), .ZN(_04799_ ) );
OAI21_X1 _19385_ ( .A(\u_lsu.pmem[1857] ), .B1(_04794_ ), .B2(_02537_ ), .ZN(_04800_ ) );
AOI21_X1 _19386_ ( .A(fanout_net_61 ), .B1(_04799_ ), .B2(_04800_ ), .ZN(_01783_ ) );
NAND3_X1 _19387_ ( .A1(_04796_ ), .A2(_03203_ ), .A3(_02535_ ), .ZN(_04801_ ) );
OAI21_X1 _19388_ ( .A(\u_lsu.pmem[1856] ), .B1(_04794_ ), .B2(_02537_ ), .ZN(_04802_ ) );
AOI21_X1 _19389_ ( .A(fanout_net_61 ), .B1(_04801_ ), .B2(_04802_ ), .ZN(_01784_ ) );
NAND4_X1 _19390_ ( .A1(_10250_ ), .A2(_04719_ ), .A3(_04732_ ), .A4(_04745_ ), .ZN(_04803_ ) );
OAI21_X1 _19391_ ( .A(\u_lsu.pmem[1831] ), .B1(_04794_ ), .B2(_02561_ ), .ZN(_04804_ ) );
AOI21_X1 _19392_ ( .A(fanout_net_61 ), .B1(_04803_ ), .B2(_04804_ ), .ZN(_01785_ ) );
BUF_X4 _19393_ ( .A(_03020_ ), .Z(_04805_ ) );
NAND4_X1 _19394_ ( .A1(_10263_ ), .A2(_04805_ ), .A3(_04732_ ), .A4(_04745_ ), .ZN(_04806_ ) );
OAI21_X1 _19395_ ( .A(\u_lsu.pmem[1830] ), .B1(_04794_ ), .B2(_02561_ ), .ZN(_04807_ ) );
AOI21_X1 _19396_ ( .A(fanout_net_61 ), .B1(_04806_ ), .B2(_04807_ ), .ZN(_01786_ ) );
NAND4_X1 _19397_ ( .A1(_10267_ ), .A2(_04805_ ), .A3(_04732_ ), .A4(_04745_ ), .ZN(_04808_ ) );
OAI21_X1 _19398_ ( .A(\u_lsu.pmem[1829] ), .B1(_04794_ ), .B2(_02561_ ), .ZN(_04809_ ) );
AOI21_X1 _19399_ ( .A(fanout_net_61 ), .B1(_04808_ ), .B2(_04809_ ), .ZN(_01787_ ) );
OAI21_X1 _19400_ ( .A(\u_lsu.pmem[4132] ), .B1(_04583_ ), .B2(_09992_ ), .ZN(_04810_ ) );
NAND4_X1 _19401_ ( .A1(_09931_ ), .A2(_04376_ ), .A3(_04556_ ), .A4(_10001_ ), .ZN(_04811_ ) );
AOI21_X1 _19402_ ( .A(fanout_net_61 ), .B1(_04810_ ), .B2(_04811_ ), .ZN(_01788_ ) );
NOR2_X1 _19403_ ( .A1(_11159_ ), .A2(_02560_ ), .ZN(_04812_ ) );
OAI21_X1 _19404_ ( .A(_09109_ ), .B1(_04812_ ), .B2(\u_lsu.pmem[1828] ), .ZN(_04813_ ) );
AOI21_X1 _19405_ ( .A(_04813_ ), .B1(_09149_ ), .B2(_04812_ ), .ZN(_01789_ ) );
NAND3_X1 _19406_ ( .A1(_04796_ ), .A2(_03114_ ), .A3(_02559_ ), .ZN(_04814_ ) );
OAI21_X1 _19407_ ( .A(\u_lsu.pmem[1827] ), .B1(_04794_ ), .B2(_02560_ ), .ZN(_04815_ ) );
AOI21_X1 _19408_ ( .A(fanout_net_61 ), .B1(_04814_ ), .B2(_04815_ ), .ZN(_01790_ ) );
NAND3_X1 _19409_ ( .A1(_04796_ ), .A2(_03145_ ), .A3(_02559_ ), .ZN(_04816_ ) );
OAI21_X1 _19410_ ( .A(\u_lsu.pmem[1826] ), .B1(_04794_ ), .B2(_02560_ ), .ZN(_04817_ ) );
AOI21_X1 _19411_ ( .A(fanout_net_62 ), .B1(_04816_ ), .B2(_04817_ ), .ZN(_01791_ ) );
NAND3_X1 _19412_ ( .A1(_04796_ ), .A2(_03174_ ), .A3(_02559_ ), .ZN(_04818_ ) );
OAI21_X1 _19413_ ( .A(\u_lsu.pmem[1825] ), .B1(_04794_ ), .B2(_02560_ ), .ZN(_04819_ ) );
AOI21_X1 _19414_ ( .A(fanout_net_62 ), .B1(_04818_ ), .B2(_04819_ ), .ZN(_01792_ ) );
BUF_X4 _19415_ ( .A(_04731_ ), .Z(_04820_ ) );
BUF_X4 _19416_ ( .A(_04685_ ), .Z(_04821_ ) );
NAND4_X1 _19417_ ( .A1(_10279_ ), .A2(_04805_ ), .A3(_04820_ ), .A4(_04821_ ), .ZN(_04822_ ) );
BUF_X4 _19418_ ( .A(_04571_ ), .Z(_04823_ ) );
OAI21_X1 _19419_ ( .A(\u_lsu.pmem[1824] ), .B1(_04823_ ), .B2(_02560_ ), .ZN(_04824_ ) );
AOI21_X1 _19420_ ( .A(fanout_net_62 ), .B1(_04822_ ), .B2(_04824_ ), .ZN(_01793_ ) );
NAND4_X1 _19421_ ( .A1(_10285_ ), .A2(_03735_ ), .A3(_04820_ ), .A4(_04821_ ), .ZN(_04825_ ) );
OAI21_X1 _19422_ ( .A(\u_lsu.pmem[1799] ), .B1(_04823_ ), .B2(_02581_ ), .ZN(_04826_ ) );
AOI21_X1 _19423_ ( .A(fanout_net_62 ), .B1(_04825_ ), .B2(_04826_ ), .ZN(_01794_ ) );
BUF_X4 _19424_ ( .A(_10287_ ), .Z(_04827_ ) );
NAND4_X1 _19425_ ( .A1(_10295_ ), .A2(_04827_ ), .A3(_04820_ ), .A4(_04821_ ), .ZN(_04828_ ) );
OAI21_X1 _19426_ ( .A(\u_lsu.pmem[1798] ), .B1(_04823_ ), .B2(_02581_ ), .ZN(_04829_ ) );
AOI21_X1 _19427_ ( .A(fanout_net_62 ), .B1(_04828_ ), .B2(_04829_ ), .ZN(_01795_ ) );
NAND4_X1 _19428_ ( .A1(_10299_ ), .A2(_04827_ ), .A3(_04820_ ), .A4(_04821_ ), .ZN(_04830_ ) );
OAI21_X1 _19429_ ( .A(\u_lsu.pmem[1797] ), .B1(_04823_ ), .B2(_02580_ ), .ZN(_04831_ ) );
AOI21_X1 _19430_ ( .A(fanout_net_62 ), .B1(_04830_ ), .B2(_04831_ ), .ZN(_01796_ ) );
NAND4_X1 _19431_ ( .A1(_10306_ ), .A2(_04827_ ), .A3(_04820_ ), .A4(_04821_ ), .ZN(_04832_ ) );
OAI21_X1 _19432_ ( .A(\u_lsu.pmem[1796] ), .B1(_04823_ ), .B2(_02580_ ), .ZN(_04833_ ) );
AOI21_X1 _19433_ ( .A(fanout_net_62 ), .B1(_04832_ ), .B2(_04833_ ), .ZN(_01797_ ) );
NAND4_X1 _19434_ ( .A1(_10309_ ), .A2(_04827_ ), .A3(_04820_ ), .A4(_04821_ ), .ZN(_04834_ ) );
OAI21_X1 _19435_ ( .A(\u_lsu.pmem[1795] ), .B1(_04823_ ), .B2(_02580_ ), .ZN(_04835_ ) );
AOI21_X1 _19436_ ( .A(fanout_net_62 ), .B1(_04834_ ), .B2(_04835_ ), .ZN(_01798_ ) );
OAI21_X1 _19437_ ( .A(\u_lsu.pmem[4131] ), .B1(_04583_ ), .B2(_09992_ ), .ZN(_04836_ ) );
NAND4_X1 _19438_ ( .A1(_03091_ ), .A2(_04376_ ), .A3(_04556_ ), .A4(_10001_ ), .ZN(_04837_ ) );
AOI21_X1 _19439_ ( .A(fanout_net_62 ), .B1(_04836_ ), .B2(_04837_ ), .ZN(_01799_ ) );
NAND4_X1 _19440_ ( .A1(_04626_ ), .A2(_04805_ ), .A3(_04820_ ), .A4(_10313_ ), .ZN(_04838_ ) );
OAI21_X1 _19441_ ( .A(\u_lsu.pmem[1794] ), .B1(_04823_ ), .B2(_02580_ ), .ZN(_04839_ ) );
AOI21_X1 _19442_ ( .A(fanout_net_62 ), .B1(_04838_ ), .B2(_04839_ ), .ZN(_01800_ ) );
NAND4_X1 _19443_ ( .A1(_10316_ ), .A2(_04827_ ), .A3(_04820_ ), .A4(_04821_ ), .ZN(_04840_ ) );
OAI21_X1 _19444_ ( .A(\u_lsu.pmem[1793] ), .B1(_04823_ ), .B2(_02580_ ), .ZN(_04841_ ) );
AOI21_X1 _19445_ ( .A(fanout_net_62 ), .B1(_04840_ ), .B2(_04841_ ), .ZN(_01801_ ) );
NAND4_X1 _19446_ ( .A1(_10320_ ), .A2(_04827_ ), .A3(_04820_ ), .A4(_04821_ ), .ZN(_04842_ ) );
OAI21_X1 _19447_ ( .A(\u_lsu.pmem[1792] ), .B1(_04823_ ), .B2(_02580_ ), .ZN(_04843_ ) );
AOI21_X1 _19448_ ( .A(fanout_net_62 ), .B1(_04842_ ), .B2(_04843_ ), .ZN(_01802_ ) );
NAND4_X1 _19449_ ( .A1(_04626_ ), .A2(_10004_ ), .A3(_09914_ ), .A4(_10324_ ), .ZN(_04844_ ) );
OAI21_X1 _19450_ ( .A(\u_lsu.pmem[1767] ), .B1(_02604_ ), .B2(_04753_ ), .ZN(_04845_ ) );
AOI21_X1 _19451_ ( .A(fanout_net_62 ), .B1(_04844_ ), .B2(_04845_ ), .ZN(_01803_ ) );
NAND4_X1 _19452_ ( .A1(_10332_ ), .A2(_04805_ ), .A3(_04820_ ), .A4(_04821_ ), .ZN(_04846_ ) );
OAI21_X1 _19453_ ( .A(\u_lsu.pmem[1766] ), .B1(_02604_ ), .B2(_04753_ ), .ZN(_04847_ ) );
AOI21_X1 _19454_ ( .A(fanout_net_62 ), .B1(_04846_ ), .B2(_04847_ ), .ZN(_01804_ ) );
BUF_X4 _19455_ ( .A(_04731_ ), .Z(_04848_ ) );
NAND4_X1 _19456_ ( .A1(_10336_ ), .A2(_04805_ ), .A3(_04848_ ), .A4(_04821_ ), .ZN(_04849_ ) );
OAI21_X1 _19457_ ( .A(\u_lsu.pmem[1765] ), .B1(_02604_ ), .B2(_04753_ ), .ZN(_04850_ ) );
AOI21_X1 _19458_ ( .A(fanout_net_62 ), .B1(_04849_ ), .B2(_04850_ ), .ZN(_01805_ ) );
BUF_X4 _19459_ ( .A(_04685_ ), .Z(_04851_ ) );
NAND4_X1 _19460_ ( .A1(_10339_ ), .A2(_04805_ ), .A3(_04848_ ), .A4(_04851_ ), .ZN(_04852_ ) );
OAI21_X1 _19461_ ( .A(\u_lsu.pmem[1764] ), .B1(_02604_ ), .B2(_04753_ ), .ZN(_04853_ ) );
AOI21_X1 _19462_ ( .A(fanout_net_62 ), .B1(_04852_ ), .B2(_04853_ ), .ZN(_01806_ ) );
NAND4_X1 _19463_ ( .A1(_10345_ ), .A2(_04805_ ), .A3(_04848_ ), .A4(_04851_ ), .ZN(_04854_ ) );
OAI21_X1 _19464_ ( .A(\u_lsu.pmem[1763] ), .B1(_02604_ ), .B2(_04753_ ), .ZN(_04855_ ) );
AOI21_X1 _19465_ ( .A(fanout_net_62 ), .B1(_04854_ ), .B2(_04855_ ), .ZN(_01807_ ) );
NAND4_X1 _19466_ ( .A1(_10350_ ), .A2(_04805_ ), .A3(_04848_ ), .A4(_04851_ ), .ZN(_04856_ ) );
OAI21_X1 _19467_ ( .A(\u_lsu.pmem[1762] ), .B1(_02604_ ), .B2(_04753_ ), .ZN(_04857_ ) );
AOI21_X1 _19468_ ( .A(fanout_net_62 ), .B1(_04856_ ), .B2(_04857_ ), .ZN(_01808_ ) );
NAND4_X1 _19469_ ( .A1(_10354_ ), .A2(_04805_ ), .A3(_04848_ ), .A4(_04851_ ), .ZN(_04858_ ) );
BUF_X4 _19470_ ( .A(_04265_ ), .Z(_04859_ ) );
OAI21_X1 _19471_ ( .A(\u_lsu.pmem[1761] ), .B1(_02604_ ), .B2(_04859_ ), .ZN(_04860_ ) );
AOI21_X1 _19472_ ( .A(fanout_net_62 ), .B1(_04858_ ), .B2(_04860_ ), .ZN(_01809_ ) );
OAI21_X1 _19473_ ( .A(\u_lsu.pmem[4130] ), .B1(_04583_ ), .B2(_09991_ ), .ZN(_04861_ ) );
BUF_X4 _19474_ ( .A(_09455_ ), .Z(_04862_ ) );
NAND4_X1 _19475_ ( .A1(_09938_ ), .A2(_04376_ ), .A3(_04862_ ), .A4(_10001_ ), .ZN(_04863_ ) );
AOI21_X1 _19476_ ( .A(fanout_net_62 ), .B1(_04861_ ), .B2(_04863_ ), .ZN(_01810_ ) );
BUF_X4 _19477_ ( .A(_03020_ ), .Z(_04864_ ) );
NAND4_X1 _19478_ ( .A1(_10357_ ), .A2(_04864_ ), .A3(_04848_ ), .A4(_04851_ ), .ZN(_04865_ ) );
OAI21_X1 _19479_ ( .A(\u_lsu.pmem[1760] ), .B1(_02604_ ), .B2(_04859_ ), .ZN(_04866_ ) );
AOI21_X1 _19480_ ( .A(fanout_net_62 ), .B1(_04865_ ), .B2(_04866_ ), .ZN(_01811_ ) );
NAND4_X1 _19481_ ( .A1(_04626_ ), .A2(_10004_ ), .A3(_09914_ ), .A4(_10362_ ), .ZN(_04867_ ) );
OAI21_X1 _19482_ ( .A(\u_lsu.pmem[1735] ), .B1(_02626_ ), .B2(_04859_ ), .ZN(_04868_ ) );
AOI21_X1 _19483_ ( .A(fanout_net_62 ), .B1(_04867_ ), .B2(_04868_ ), .ZN(_01812_ ) );
NAND4_X1 _19484_ ( .A1(_10368_ ), .A2(_04864_ ), .A3(_04848_ ), .A4(_04851_ ), .ZN(_04869_ ) );
OAI21_X1 _19485_ ( .A(\u_lsu.pmem[1734] ), .B1(_02626_ ), .B2(_04859_ ), .ZN(_04870_ ) );
AOI21_X1 _19486_ ( .A(fanout_net_62 ), .B1(_04869_ ), .B2(_04870_ ), .ZN(_01813_ ) );
NAND4_X1 _19487_ ( .A1(_10371_ ), .A2(_04864_ ), .A3(_04848_ ), .A4(_04851_ ), .ZN(_04871_ ) );
OAI21_X1 _19488_ ( .A(\u_lsu.pmem[1733] ), .B1(_02626_ ), .B2(_04859_ ), .ZN(_04872_ ) );
AOI21_X1 _19489_ ( .A(fanout_net_62 ), .B1(_04871_ ), .B2(_04872_ ), .ZN(_01814_ ) );
NAND4_X1 _19490_ ( .A1(_10374_ ), .A2(_04864_ ), .A3(_04848_ ), .A4(_04851_ ), .ZN(_04873_ ) );
OAI21_X1 _19491_ ( .A(\u_lsu.pmem[1732] ), .B1(_02626_ ), .B2(_04859_ ), .ZN(_04874_ ) );
AOI21_X1 _19492_ ( .A(fanout_net_62 ), .B1(_04873_ ), .B2(_04874_ ), .ZN(_01815_ ) );
NAND4_X1 _19493_ ( .A1(_10377_ ), .A2(_04864_ ), .A3(_04848_ ), .A4(_04851_ ), .ZN(_04875_ ) );
OAI21_X1 _19494_ ( .A(\u_lsu.pmem[1731] ), .B1(_02626_ ), .B2(_04859_ ), .ZN(_04876_ ) );
AOI21_X1 _19495_ ( .A(fanout_net_62 ), .B1(_04875_ ), .B2(_04876_ ), .ZN(_01816_ ) );
BUF_X4 _19496_ ( .A(_04731_ ), .Z(_04877_ ) );
NAND4_X1 _19497_ ( .A1(_10381_ ), .A2(_04864_ ), .A3(_04877_ ), .A4(_04851_ ), .ZN(_04878_ ) );
OAI21_X1 _19498_ ( .A(\u_lsu.pmem[1730] ), .B1(_02626_ ), .B2(_04859_ ), .ZN(_04879_ ) );
AOI21_X1 _19499_ ( .A(fanout_net_62 ), .B1(_04878_ ), .B2(_04879_ ), .ZN(_01817_ ) );
BUF_X4 _19500_ ( .A(_04685_ ), .Z(_04880_ ) );
NAND4_X1 _19501_ ( .A1(_10384_ ), .A2(_04864_ ), .A3(_04877_ ), .A4(_04880_ ), .ZN(_04881_ ) );
OAI21_X1 _19502_ ( .A(\u_lsu.pmem[1729] ), .B1(_02626_ ), .B2(_04859_ ), .ZN(_04882_ ) );
AOI21_X1 _19503_ ( .A(fanout_net_62 ), .B1(_04881_ ), .B2(_04882_ ), .ZN(_01818_ ) );
NAND4_X1 _19504_ ( .A1(_10391_ ), .A2(_04864_ ), .A3(_04877_ ), .A4(_04880_ ), .ZN(_04883_ ) );
OAI21_X1 _19505_ ( .A(\u_lsu.pmem[1728] ), .B1(_02626_ ), .B2(_04859_ ), .ZN(_04884_ ) );
AOI21_X1 _19506_ ( .A(fanout_net_62 ), .B1(_04883_ ), .B2(_04884_ ), .ZN(_01819_ ) );
NAND4_X1 _19507_ ( .A1(_10394_ ), .A2(_04864_ ), .A3(_04877_ ), .A4(_04880_ ), .ZN(_04885_ ) );
BUF_X4 _19508_ ( .A(_04265_ ), .Z(_04886_ ) );
OAI21_X1 _19509_ ( .A(\u_lsu.pmem[1703] ), .B1(_02650_ ), .B2(_04886_ ), .ZN(_04887_ ) );
AOI21_X1 _19510_ ( .A(fanout_net_62 ), .B1(_04885_ ), .B2(_04887_ ), .ZN(_01820_ ) );
OAI21_X1 _19511_ ( .A(\u_lsu.pmem[4129] ), .B1(_04583_ ), .B2(_09991_ ), .ZN(_04888_ ) );
NAND4_X1 _19512_ ( .A1(_03143_ ), .A2(_04376_ ), .A3(_04862_ ), .A4(_09990_ ), .ZN(_04889_ ) );
AOI21_X1 _19513_ ( .A(fanout_net_63 ), .B1(_04888_ ), .B2(_04889_ ), .ZN(_01821_ ) );
NAND4_X1 _19514_ ( .A1(_10402_ ), .A2(_04864_ ), .A3(_04877_ ), .A4(_04880_ ), .ZN(_04890_ ) );
OAI21_X1 _19515_ ( .A(\u_lsu.pmem[1702] ), .B1(_02650_ ), .B2(_04886_ ), .ZN(_04891_ ) );
AOI21_X1 _19516_ ( .A(fanout_net_63 ), .B1(_04890_ ), .B2(_04891_ ), .ZN(_01822_ ) );
BUF_X4 _19517_ ( .A(_03020_ ), .Z(_04892_ ) );
NAND4_X1 _19518_ ( .A1(_10405_ ), .A2(_04892_ ), .A3(_04877_ ), .A4(_04880_ ), .ZN(_04893_ ) );
OAI21_X1 _19519_ ( .A(\u_lsu.pmem[1701] ), .B1(_02650_ ), .B2(_04886_ ), .ZN(_04894_ ) );
AOI21_X1 _19520_ ( .A(fanout_net_63 ), .B1(_04893_ ), .B2(_04894_ ), .ZN(_01823_ ) );
NAND4_X1 _19521_ ( .A1(_10408_ ), .A2(_04892_ ), .A3(_04877_ ), .A4(_04880_ ), .ZN(_04895_ ) );
OAI21_X1 _19522_ ( .A(\u_lsu.pmem[1700] ), .B1(_02650_ ), .B2(_04886_ ), .ZN(_04896_ ) );
AOI21_X1 _19523_ ( .A(fanout_net_63 ), .B1(_04895_ ), .B2(_04896_ ), .ZN(_01824_ ) );
NAND4_X1 _19524_ ( .A1(_10411_ ), .A2(_04892_ ), .A3(_04877_ ), .A4(_04880_ ), .ZN(_04897_ ) );
OAI21_X1 _19525_ ( .A(\u_lsu.pmem[1699] ), .B1(_02650_ ), .B2(_04886_ ), .ZN(_04898_ ) );
AOI21_X1 _19526_ ( .A(fanout_net_63 ), .B1(_04897_ ), .B2(_04898_ ), .ZN(_01825_ ) );
NAND4_X1 _19527_ ( .A1(_10414_ ), .A2(_04892_ ), .A3(_04877_ ), .A4(_04880_ ), .ZN(_04899_ ) );
OAI21_X1 _19528_ ( .A(\u_lsu.pmem[1698] ), .B1(_02650_ ), .B2(_04886_ ), .ZN(_04900_ ) );
AOI21_X1 _19529_ ( .A(fanout_net_63 ), .B1(_04899_ ), .B2(_04900_ ), .ZN(_01826_ ) );
NAND4_X1 _19530_ ( .A1(_10417_ ), .A2(_04892_ ), .A3(_04877_ ), .A4(_04880_ ), .ZN(_04901_ ) );
OAI21_X1 _19531_ ( .A(\u_lsu.pmem[1697] ), .B1(_02650_ ), .B2(_04886_ ), .ZN(_04902_ ) );
AOI21_X1 _19532_ ( .A(fanout_net_63 ), .B1(_04901_ ), .B2(_04902_ ), .ZN(_01827_ ) );
BUF_X4 _19533_ ( .A(_09953_ ), .Z(_04903_ ) );
NAND4_X1 _19534_ ( .A1(_04903_ ), .A2(_10004_ ), .A3(_03753_ ), .A4(_10398_ ), .ZN(_04904_ ) );
OAI21_X1 _19535_ ( .A(\u_lsu.pmem[1696] ), .B1(_02650_ ), .B2(_04886_ ), .ZN(_04905_ ) );
AOI21_X1 _19536_ ( .A(fanout_net_63 ), .B1(_04904_ ), .B2(_04905_ ), .ZN(_01828_ ) );
OAI21_X1 _19537_ ( .A(\u_lsu.pmem[1671] ), .B1(_02678_ ), .B2(_04593_ ), .ZN(_04906_ ) );
NAND4_X1 _19538_ ( .A1(_10436_ ), .A2(_03107_ ), .A3(_04862_ ), .A4(_04595_ ), .ZN(_04907_ ) );
AOI21_X1 _19539_ ( .A(fanout_net_63 ), .B1(_04906_ ), .B2(_04907_ ), .ZN(_01829_ ) );
BUF_X4 _19540_ ( .A(_04731_ ), .Z(_04908_ ) );
NAND4_X1 _19541_ ( .A1(_02682_ ), .A2(_09658_ ), .A3(_04908_ ), .A4(_04880_ ), .ZN(_04909_ ) );
OAI21_X1 _19542_ ( .A(\u_lsu.pmem[1670] ), .B1(_02677_ ), .B2(_04886_ ), .ZN(_04910_ ) );
AOI21_X1 _19543_ ( .A(fanout_net_63 ), .B1(_04909_ ), .B2(_04910_ ), .ZN(_01830_ ) );
BUF_X4 _19544_ ( .A(_04685_ ), .Z(_04911_ ) );
NAND4_X1 _19545_ ( .A1(_02682_ ), .A2(_09713_ ), .A3(_04908_ ), .A4(_04911_ ), .ZN(_04912_ ) );
OAI21_X1 _19546_ ( .A(\u_lsu.pmem[1669] ), .B1(_02677_ ), .B2(_04886_ ), .ZN(_04913_ ) );
AOI21_X1 _19547_ ( .A(fanout_net_63 ), .B1(_04912_ ), .B2(_04913_ ), .ZN(_01831_ ) );
BUF_X4 _19548_ ( .A(_04210_ ), .Z(_04914_ ) );
NAND4_X1 _19549_ ( .A1(_10021_ ), .A2(_04914_ ), .A3(_04908_ ), .A4(_04097_ ), .ZN(_04915_ ) );
OAI21_X1 _19550_ ( .A(\u_lsu.pmem[4128] ), .B1(_04071_ ), .B2(_09991_ ), .ZN(_04916_ ) );
AOI21_X1 _19551_ ( .A(fanout_net_63 ), .B1(_04915_ ), .B2(_04916_ ), .ZN(_01832_ ) );
NAND4_X1 _19552_ ( .A1(_10442_ ), .A2(_09514_ ), .A3(_04908_ ), .A4(_04911_ ), .ZN(_04917_ ) );
BUF_X4 _19553_ ( .A(_04265_ ), .Z(_04918_ ) );
OAI21_X1 _19554_ ( .A(\u_lsu.pmem[1668] ), .B1(_02677_ ), .B2(_04918_ ), .ZN(_04919_ ) );
AOI21_X1 _19555_ ( .A(fanout_net_63 ), .B1(_04917_ ), .B2(_04919_ ), .ZN(_01833_ ) );
NAND4_X1 _19556_ ( .A1(_10442_ ), .A2(_09520_ ), .A3(_04908_ ), .A4(_04911_ ), .ZN(_04920_ ) );
OAI21_X1 _19557_ ( .A(\u_lsu.pmem[1667] ), .B1(_02677_ ), .B2(_04918_ ), .ZN(_04921_ ) );
AOI21_X1 _19558_ ( .A(fanout_net_63 ), .B1(_04920_ ), .B2(_04921_ ), .ZN(_01834_ ) );
OAI21_X1 _19559_ ( .A(\u_lsu.pmem[1666] ), .B1(_02678_ ), .B2(_04593_ ), .ZN(_04922_ ) );
NAND4_X1 _19560_ ( .A1(_10460_ ), .A2(_10126_ ), .A3(_04862_ ), .A4(_04595_ ), .ZN(_04923_ ) );
AOI21_X1 _19561_ ( .A(fanout_net_63 ), .B1(_04922_ ), .B2(_04923_ ), .ZN(_01835_ ) );
NAND4_X1 _19562_ ( .A1(_10442_ ), .A2(_09544_ ), .A3(_04908_ ), .A4(_04911_ ), .ZN(_04924_ ) );
OAI21_X1 _19563_ ( .A(\u_lsu.pmem[1665] ), .B1(_02677_ ), .B2(_04918_ ), .ZN(_04925_ ) );
AOI21_X1 _19564_ ( .A(fanout_net_63 ), .B1(_04924_ ), .B2(_04925_ ), .ZN(_01836_ ) );
NAND4_X1 _19565_ ( .A1(_10442_ ), .A2(_09548_ ), .A3(_04908_ ), .A4(_04911_ ), .ZN(_04926_ ) );
OAI21_X1 _19566_ ( .A(\u_lsu.pmem[1664] ), .B1(_02677_ ), .B2(_04918_ ), .ZN(_04927_ ) );
AOI21_X1 _19567_ ( .A(fanout_net_63 ), .B1(_04926_ ), .B2(_04927_ ), .ZN(_01837_ ) );
BUF_X4 _19568_ ( .A(_09566_ ), .Z(_04928_ ) );
NAND4_X1 _19569_ ( .A1(_04903_ ), .A2(_10004_ ), .A3(_04928_ ), .A4(_02757_ ), .ZN(_04929_ ) );
OAI21_X1 _19570_ ( .A(\u_lsu.pmem[1639] ), .B1(_02700_ ), .B2(_04918_ ), .ZN(_04930_ ) );
AOI21_X1 _19571_ ( .A(fanout_net_63 ), .B1(_04929_ ), .B2(_04930_ ), .ZN(_01838_ ) );
NAND4_X1 _19572_ ( .A1(_04903_ ), .A2(_10004_ ), .A3(_09925_ ), .A4(_02757_ ), .ZN(_04931_ ) );
OAI21_X1 _19573_ ( .A(\u_lsu.pmem[1638] ), .B1(_02700_ ), .B2(_04918_ ), .ZN(_04932_ ) );
AOI21_X1 _19574_ ( .A(fanout_net_63 ), .B1(_04931_ ), .B2(_04932_ ), .ZN(_01839_ ) );
NAND4_X1 _19575_ ( .A1(_04903_ ), .A2(_10004_ ), .A3(_09928_ ), .A4(_10475_ ), .ZN(_04933_ ) );
OAI21_X1 _19576_ ( .A(\u_lsu.pmem[1637] ), .B1(_02700_ ), .B2(_04918_ ), .ZN(_04934_ ) );
AOI21_X1 _19577_ ( .A(fanout_net_63 ), .B1(_04933_ ), .B2(_04934_ ), .ZN(_01840_ ) );
NAND4_X1 _19578_ ( .A1(_04903_ ), .A2(_10004_ ), .A3(_11151_ ), .A4(_10475_ ), .ZN(_04935_ ) );
OAI21_X1 _19579_ ( .A(\u_lsu.pmem[1636] ), .B1(_02700_ ), .B2(_04918_ ), .ZN(_04936_ ) );
AOI21_X1 _19580_ ( .A(fanout_net_63 ), .B1(_04935_ ), .B2(_04936_ ), .ZN(_01841_ ) );
BUF_X4 _19581_ ( .A(_09456_ ), .Z(_04937_ ) );
NAND4_X1 _19582_ ( .A1(_04903_ ), .A2(_04937_ ), .A3(_09934_ ), .A4(_10475_ ), .ZN(_04938_ ) );
OAI21_X1 _19583_ ( .A(\u_lsu.pmem[1635] ), .B1(_02700_ ), .B2(_04918_ ), .ZN(_04939_ ) );
AOI21_X1 _19584_ ( .A(fanout_net_63 ), .B1(_04938_ ), .B2(_04939_ ), .ZN(_01842_ ) );
AND2_X1 _19585_ ( .A1(_09498_ ), .A2(_10045_ ), .ZN(_04940_ ) );
INV_X1 _19586_ ( .A(_04940_ ), .ZN(_04941_ ) );
NAND2_X1 _19587_ ( .A1(_04941_ ), .A2(\u_lsu.pmem[4103] ), .ZN(_04942_ ) );
NAND4_X1 _19588_ ( .A1(_04669_ ), .A2(_03478_ ), .A3(_10589_ ), .A4(_02485_ ), .ZN(_04943_ ) );
AOI21_X1 _19589_ ( .A(fanout_net_63 ), .B1(_04942_ ), .B2(_04943_ ), .ZN(_01843_ ) );
NAND4_X1 _19590_ ( .A1(_04903_ ), .A2(_04937_ ), .A3(_10015_ ), .A4(_10475_ ), .ZN(_04944_ ) );
OAI21_X1 _19591_ ( .A(\u_lsu.pmem[1634] ), .B1(_02700_ ), .B2(_04918_ ), .ZN(_04945_ ) );
AOI21_X1 _19592_ ( .A(fanout_net_63 ), .B1(_04944_ ), .B2(_04945_ ), .ZN(_01844_ ) );
NAND4_X1 _19593_ ( .A1(_04903_ ), .A2(_04937_ ), .A3(_09941_ ), .A4(_10475_ ), .ZN(_04946_ ) );
BUF_X4 _19594_ ( .A(_04265_ ), .Z(_04947_ ) );
OAI21_X1 _19595_ ( .A(\u_lsu.pmem[1633] ), .B1(_02700_ ), .B2(_04947_ ), .ZN(_04948_ ) );
AOI21_X1 _19596_ ( .A(fanout_net_63 ), .B1(_04946_ ), .B2(_04948_ ), .ZN(_01845_ ) );
NAND4_X1 _19597_ ( .A1(_04903_ ), .A2(_04937_ ), .A3(_03753_ ), .A4(_10475_ ), .ZN(_04949_ ) );
OAI21_X1 _19598_ ( .A(\u_lsu.pmem[1632] ), .B1(_02700_ ), .B2(_04947_ ), .ZN(_04950_ ) );
AOI21_X1 _19599_ ( .A(fanout_net_63 ), .B1(_04949_ ), .B2(_04950_ ), .ZN(_01846_ ) );
NAND4_X1 _19600_ ( .A1(_04903_ ), .A2(_04937_ ), .A3(_04928_ ), .A4(_10506_ ), .ZN(_04951_ ) );
OAI21_X1 _19601_ ( .A(\u_lsu.pmem[1607] ), .B1(_02723_ ), .B2(_04947_ ), .ZN(_04952_ ) );
AOI21_X1 _19602_ ( .A(fanout_net_63 ), .B1(_04951_ ), .B2(_04952_ ), .ZN(_01847_ ) );
BUF_X4 _19603_ ( .A(_09953_ ), .Z(_04953_ ) );
NAND4_X1 _19604_ ( .A1(_04953_ ), .A2(_04937_ ), .A3(_09925_ ), .A4(_10506_ ), .ZN(_04954_ ) );
OAI21_X1 _19605_ ( .A(\u_lsu.pmem[1606] ), .B1(_02723_ ), .B2(_04947_ ), .ZN(_04955_ ) );
AOI21_X1 _19606_ ( .A(fanout_net_63 ), .B1(_04954_ ), .B2(_04955_ ), .ZN(_01848_ ) );
NAND4_X1 _19607_ ( .A1(_04953_ ), .A2(_04937_ ), .A3(_09928_ ), .A4(_10506_ ), .ZN(_04956_ ) );
OAI21_X1 _19608_ ( .A(\u_lsu.pmem[1605] ), .B1(_02723_ ), .B2(_04947_ ), .ZN(_04957_ ) );
AOI21_X1 _19609_ ( .A(fanout_net_63 ), .B1(_04956_ ), .B2(_04957_ ), .ZN(_01849_ ) );
NAND4_X1 _19610_ ( .A1(_04953_ ), .A2(_04937_ ), .A3(_11151_ ), .A4(_10506_ ), .ZN(_04958_ ) );
OAI21_X1 _19611_ ( .A(\u_lsu.pmem[1604] ), .B1(_02723_ ), .B2(_04947_ ), .ZN(_04959_ ) );
AOI21_X1 _19612_ ( .A(fanout_net_63 ), .B1(_04958_ ), .B2(_04959_ ), .ZN(_01850_ ) );
NAND4_X1 _19613_ ( .A1(_04953_ ), .A2(_04937_ ), .A3(_09934_ ), .A4(_10506_ ), .ZN(_04960_ ) );
OAI21_X1 _19614_ ( .A(\u_lsu.pmem[1603] ), .B1(_02723_ ), .B2(_04947_ ), .ZN(_04961_ ) );
AOI21_X1 _19615_ ( .A(fanout_net_64 ), .B1(_04960_ ), .B2(_04961_ ), .ZN(_01851_ ) );
NAND4_X1 _19616_ ( .A1(_04953_ ), .A2(_04937_ ), .A3(_10015_ ), .A4(_10506_ ), .ZN(_04962_ ) );
OAI21_X1 _19617_ ( .A(\u_lsu.pmem[1602] ), .B1(_02723_ ), .B2(_04947_ ), .ZN(_04963_ ) );
AOI21_X1 _19618_ ( .A(fanout_net_64 ), .B1(_04962_ ), .B2(_04963_ ), .ZN(_01852_ ) );
BUF_X4 _19619_ ( .A(_09456_ ), .Z(_04964_ ) );
NAND4_X1 _19620_ ( .A1(_04953_ ), .A2(_04964_ ), .A3(_09941_ ), .A4(_10506_ ), .ZN(_04965_ ) );
OAI21_X1 _19621_ ( .A(\u_lsu.pmem[1601] ), .B1(_02723_ ), .B2(_04947_ ), .ZN(_04966_ ) );
AOI21_X1 _19622_ ( .A(fanout_net_64 ), .B1(_04965_ ), .B2(_04966_ ), .ZN(_01853_ ) );
NAND4_X1 _19623_ ( .A1(_09718_ ), .A2(_04914_ ), .A3(_04908_ ), .A4(_04097_ ), .ZN(_04967_ ) );
OAI21_X1 _19624_ ( .A(\u_lsu.pmem[4357] ), .B1(_04071_ ), .B2(_09468_ ), .ZN(_04968_ ) );
AOI21_X1 _19625_ ( .A(fanout_net_64 ), .B1(_04967_ ), .B2(_04968_ ), .ZN(_01854_ ) );
NAND2_X1 _19626_ ( .A1(_04941_ ), .A2(\u_lsu.pmem[4102] ), .ZN(_04969_ ) );
NAND4_X1 _19627_ ( .A1(_04669_ ), .A2(_09575_ ), .A3(_10589_ ), .A4(_02485_ ), .ZN(_04970_ ) );
AOI21_X1 _19628_ ( .A(fanout_net_64 ), .B1(_04969_ ), .B2(_04970_ ), .ZN(_01855_ ) );
NAND4_X1 _19629_ ( .A1(_04953_ ), .A2(_04964_ ), .A3(_03753_ ), .A4(_10506_ ), .ZN(_04971_ ) );
OAI21_X1 _19630_ ( .A(\u_lsu.pmem[1600] ), .B1(_02723_ ), .B2(_04947_ ), .ZN(_04972_ ) );
AOI21_X1 _19631_ ( .A(fanout_net_64 ), .B1(_04971_ ), .B2(_04972_ ), .ZN(_01856_ ) );
NAND4_X1 _19632_ ( .A1(_10527_ ), .A2(_04892_ ), .A3(_04908_ ), .A4(_04911_ ), .ZN(_04973_ ) );
BUF_X4 _19633_ ( .A(_04265_ ), .Z(_04974_ ) );
OAI21_X1 _19634_ ( .A(\u_lsu.pmem[1575] ), .B1(_02751_ ), .B2(_04974_ ), .ZN(_04975_ ) );
AOI21_X1 _19635_ ( .A(fanout_net_64 ), .B1(_04973_ ), .B2(_04975_ ), .ZN(_01857_ ) );
NAND4_X1 _19636_ ( .A1(_10535_ ), .A2(_04892_ ), .A3(_04908_ ), .A4(_04911_ ), .ZN(_04976_ ) );
OAI21_X1 _19637_ ( .A(\u_lsu.pmem[1574] ), .B1(_02751_ ), .B2(_04974_ ), .ZN(_04977_ ) );
AOI21_X1 _19638_ ( .A(fanout_net_64 ), .B1(_04976_ ), .B2(_04977_ ), .ZN(_01858_ ) );
BUF_X4 _19639_ ( .A(_04731_ ), .Z(_04978_ ) );
NAND4_X1 _19640_ ( .A1(_10538_ ), .A2(_04892_ ), .A3(_04978_ ), .A4(_04911_ ), .ZN(_04979_ ) );
OAI21_X1 _19641_ ( .A(\u_lsu.pmem[1573] ), .B1(_02751_ ), .B2(_04974_ ), .ZN(_04980_ ) );
AOI21_X1 _19642_ ( .A(fanout_net_64 ), .B1(_04979_ ), .B2(_04980_ ), .ZN(_01859_ ) );
NAND4_X1 _19643_ ( .A1(_04953_ ), .A2(_04964_ ), .A3(_11151_ ), .A4(_10542_ ), .ZN(_04981_ ) );
OAI21_X1 _19644_ ( .A(\u_lsu.pmem[1572] ), .B1(_02751_ ), .B2(_04974_ ), .ZN(_04982_ ) );
AOI21_X1 _19645_ ( .A(fanout_net_64 ), .B1(_04981_ ), .B2(_04982_ ), .ZN(_01860_ ) );
NAND4_X1 _19646_ ( .A1(_04953_ ), .A2(_04964_ ), .A3(_09934_ ), .A4(_10542_ ), .ZN(_04983_ ) );
OAI21_X1 _19647_ ( .A(\u_lsu.pmem[1571] ), .B1(_02751_ ), .B2(_04974_ ), .ZN(_04984_ ) );
AOI21_X1 _19648_ ( .A(fanout_net_64 ), .B1(_04983_ ), .B2(_04984_ ), .ZN(_01861_ ) );
NAND4_X1 _19649_ ( .A1(_04953_ ), .A2(_04964_ ), .A3(_10015_ ), .A4(_10542_ ), .ZN(_04985_ ) );
OAI21_X1 _19650_ ( .A(\u_lsu.pmem[1570] ), .B1(_02751_ ), .B2(_04974_ ), .ZN(_04986_ ) );
AOI21_X1 _19651_ ( .A(fanout_net_64 ), .B1(_04985_ ), .B2(_04986_ ), .ZN(_01862_ ) );
BUF_X4 _19652_ ( .A(_09953_ ), .Z(_04987_ ) );
NAND4_X1 _19653_ ( .A1(_04987_ ), .A2(_04964_ ), .A3(_09941_ ), .A4(_10542_ ), .ZN(_04988_ ) );
OAI21_X1 _19654_ ( .A(\u_lsu.pmem[1569] ), .B1(_02751_ ), .B2(_04974_ ), .ZN(_04989_ ) );
AOI21_X1 _19655_ ( .A(fanout_net_64 ), .B1(_04988_ ), .B2(_04989_ ), .ZN(_01863_ ) );
NAND4_X1 _19656_ ( .A1(_10556_ ), .A2(_04892_ ), .A3(_04978_ ), .A4(_04911_ ), .ZN(_04990_ ) );
OAI21_X1 _19657_ ( .A(\u_lsu.pmem[1568] ), .B1(_02751_ ), .B2(_04974_ ), .ZN(_04991_ ) );
AOI21_X1 _19658_ ( .A(fanout_net_64 ), .B1(_04990_ ), .B2(_04991_ ), .ZN(_01864_ ) );
NAND3_X1 _19659_ ( .A1(_04796_ ), .A2(_11423_ ), .A3(_02772_ ), .ZN(_04992_ ) );
OAI21_X1 _19660_ ( .A(\u_lsu.pmem[1543] ), .B1(_04823_ ), .B2(_02770_ ), .ZN(_04993_ ) );
AOI21_X1 _19661_ ( .A(fanout_net_64 ), .B1(_04992_ ), .B2(_04993_ ), .ZN(_01865_ ) );
NAND2_X1 _19662_ ( .A1(_04941_ ), .A2(\u_lsu.pmem[4101] ), .ZN(_04994_ ) );
NAND4_X1 _19663_ ( .A1(_04669_ ), .A2(_09582_ ), .A3(_10589_ ), .A4(_02485_ ), .ZN(_04995_ ) );
AOI21_X1 _19664_ ( .A(fanout_net_64 ), .B1(_04994_ ), .B2(_04995_ ), .ZN(_01866_ ) );
NAND3_X1 _19665_ ( .A1(_04796_ ), .A2(_10444_ ), .A3(_02772_ ), .ZN(_04996_ ) );
BUF_X4 _19666_ ( .A(_04571_ ), .Z(_04997_ ) );
OAI21_X1 _19667_ ( .A(\u_lsu.pmem[1542] ), .B1(_04997_ ), .B2(_02770_ ), .ZN(_04998_ ) );
AOI21_X1 _19668_ ( .A(fanout_net_64 ), .B1(_04996_ ), .B2(_04998_ ), .ZN(_01867_ ) );
NAND3_X1 _19669_ ( .A1(_04796_ ), .A2(_10448_ ), .A3(_02772_ ), .ZN(_04999_ ) );
OAI21_X1 _19670_ ( .A(\u_lsu.pmem[1541] ), .B1(_04997_ ), .B2(_02769_ ), .ZN(_05000_ ) );
AOI21_X1 _19671_ ( .A(fanout_net_64 ), .B1(_04999_ ), .B2(_05000_ ), .ZN(_01868_ ) );
NAND3_X1 _19672_ ( .A1(_04796_ ), .A2(_10453_ ), .A3(_02772_ ), .ZN(_05001_ ) );
OAI21_X1 _19673_ ( .A(\u_lsu.pmem[1540] ), .B1(_04997_ ), .B2(_02769_ ), .ZN(_05002_ ) );
AOI21_X1 _19674_ ( .A(fanout_net_64 ), .B1(_05001_ ), .B2(_05002_ ), .ZN(_01869_ ) );
NAND4_X1 _19675_ ( .A1(_10575_ ), .A2(_04827_ ), .A3(_04978_ ), .A4(_04911_ ), .ZN(_05003_ ) );
OAI21_X1 _19676_ ( .A(\u_lsu.pmem[1539] ), .B1(_04997_ ), .B2(_02769_ ), .ZN(_05004_ ) );
AOI21_X1 _19677_ ( .A(fanout_net_64 ), .B1(_05003_ ), .B2(_05004_ ), .ZN(_01870_ ) );
BUF_X4 _19678_ ( .A(_04685_ ), .Z(_05005_ ) );
NAND4_X1 _19679_ ( .A1(_10584_ ), .A2(_02486_ ), .A3(_10876_ ), .A4(_05005_ ), .ZN(_05006_ ) );
OAI21_X1 _19680_ ( .A(\u_lsu.pmem[1538] ), .B1(_04997_ ), .B2(_02769_ ), .ZN(_05007_ ) );
AOI21_X1 _19681_ ( .A(fanout_net_64 ), .B1(_05006_ ), .B2(_05007_ ), .ZN(_01871_ ) );
BUF_X4 _19682_ ( .A(_09641_ ), .Z(_05008_ ) );
NAND3_X1 _19683_ ( .A1(_05008_ ), .A2(_10463_ ), .A3(_02772_ ), .ZN(_05009_ ) );
OAI21_X1 _19684_ ( .A(\u_lsu.pmem[1537] ), .B1(_04997_ ), .B2(_02769_ ), .ZN(_05010_ ) );
AOI21_X1 _19685_ ( .A(fanout_net_64 ), .B1(_05009_ ), .B2(_05010_ ), .ZN(_01872_ ) );
BUF_X4 _19686_ ( .A(_09476_ ), .Z(_05011_ ) );
NAND4_X1 _19687_ ( .A1(_10591_ ), .A2(_09676_ ), .A3(_03673_ ), .A4(_05011_ ), .ZN(_05012_ ) );
OAI21_X1 _19688_ ( .A(\u_lsu.pmem[1536] ), .B1(_04997_ ), .B2(_02769_ ), .ZN(_05013_ ) );
AOI21_X1 _19689_ ( .A(fanout_net_64 ), .B1(_05012_ ), .B2(_05013_ ), .ZN(_01873_ ) );
NAND4_X1 _19690_ ( .A1(_04987_ ), .A2(_04964_ ), .A3(_04928_ ), .A4(_10596_ ), .ZN(_05014_ ) );
OAI21_X1 _19691_ ( .A(\u_lsu.pmem[1511] ), .B1(_02793_ ), .B2(_04974_ ), .ZN(_05015_ ) );
AOI21_X1 _19692_ ( .A(fanout_net_64 ), .B1(_05014_ ), .B2(_05015_ ), .ZN(_01874_ ) );
NAND4_X1 _19693_ ( .A1(_10603_ ), .A2(_04892_ ), .A3(_04978_ ), .A4(_05005_ ), .ZN(_05016_ ) );
OAI21_X1 _19694_ ( .A(\u_lsu.pmem[1510] ), .B1(_02793_ ), .B2(_04974_ ), .ZN(_05017_ ) );
AOI21_X1 _19695_ ( .A(fanout_net_64 ), .B1(_05016_ ), .B2(_05017_ ), .ZN(_01875_ ) );
NAND4_X1 _19696_ ( .A1(_10608_ ), .A2(_04827_ ), .A3(_04978_ ), .A4(_05005_ ), .ZN(_05018_ ) );
BUF_X4 _19697_ ( .A(_04265_ ), .Z(_05019_ ) );
OAI21_X1 _19698_ ( .A(\u_lsu.pmem[1509] ), .B1(_02793_ ), .B2(_05019_ ), .ZN(_05020_ ) );
AOI21_X1 _19699_ ( .A(fanout_net_64 ), .B1(_05018_ ), .B2(_05020_ ), .ZN(_01876_ ) );
NAND2_X1 _19700_ ( .A1(_04941_ ), .A2(\u_lsu.pmem[4100] ), .ZN(_05021_ ) );
NAND4_X1 _19701_ ( .A1(_04669_ ), .A2(_08605_ ), .A3(_10589_ ), .A4(_02485_ ), .ZN(_05022_ ) );
AOI21_X1 _19702_ ( .A(fanout_net_64 ), .B1(_05021_ ), .B2(_05022_ ), .ZN(_01877_ ) );
NAND4_X1 _19703_ ( .A1(_10611_ ), .A2(_04827_ ), .A3(_04978_ ), .A4(_05005_ ), .ZN(_05023_ ) );
OAI21_X1 _19704_ ( .A(\u_lsu.pmem[1508] ), .B1(_02793_ ), .B2(_05019_ ), .ZN(_05024_ ) );
AOI21_X1 _19705_ ( .A(fanout_net_64 ), .B1(_05023_ ), .B2(_05024_ ), .ZN(_01878_ ) );
NAND4_X1 _19706_ ( .A1(_10614_ ), .A2(_04827_ ), .A3(_04978_ ), .A4(_05005_ ), .ZN(_05025_ ) );
OAI21_X1 _19707_ ( .A(\u_lsu.pmem[1507] ), .B1(_02793_ ), .B2(_05019_ ), .ZN(_05026_ ) );
AOI21_X1 _19708_ ( .A(fanout_net_64 ), .B1(_05025_ ), .B2(_05026_ ), .ZN(_01879_ ) );
BUF_X4 _19709_ ( .A(_10287_ ), .Z(_05027_ ) );
NAND4_X1 _19710_ ( .A1(_10617_ ), .A2(_05027_ ), .A3(_04978_ ), .A4(_05005_ ), .ZN(_05028_ ) );
OAI21_X1 _19711_ ( .A(\u_lsu.pmem[1506] ), .B1(_02793_ ), .B2(_05019_ ), .ZN(_05029_ ) );
AOI21_X1 _19712_ ( .A(fanout_net_64 ), .B1(_05028_ ), .B2(_05029_ ), .ZN(_01880_ ) );
BUF_X4 _19713_ ( .A(_10063_ ), .Z(_05030_ ) );
NAND4_X1 _19714_ ( .A1(_10621_ ), .A2(_05030_ ), .A3(_04978_ ), .A4(_05005_ ), .ZN(_05031_ ) );
OAI21_X1 _19715_ ( .A(\u_lsu.pmem[1505] ), .B1(_02793_ ), .B2(_05019_ ), .ZN(_05032_ ) );
AOI21_X1 _19716_ ( .A(fanout_net_65 ), .B1(_05031_ ), .B2(_05032_ ), .ZN(_01881_ ) );
NAND4_X1 _19717_ ( .A1(_10624_ ), .A2(_05027_ ), .A3(_04978_ ), .A4(_05005_ ), .ZN(_05033_ ) );
OAI21_X1 _19718_ ( .A(\u_lsu.pmem[1504] ), .B1(_02793_ ), .B2(_05019_ ), .ZN(_05034_ ) );
AOI21_X1 _19719_ ( .A(fanout_net_65 ), .B1(_05033_ ), .B2(_05034_ ), .ZN(_01882_ ) );
NAND4_X1 _19720_ ( .A1(_04987_ ), .A2(_04964_ ), .A3(_04928_ ), .A4(_10627_ ), .ZN(_05035_ ) );
OAI21_X1 _19721_ ( .A(\u_lsu.pmem[1479] ), .B1(_02814_ ), .B2(_05019_ ), .ZN(_05036_ ) );
AOI21_X1 _19722_ ( .A(fanout_net_65 ), .B1(_05035_ ), .B2(_05036_ ), .ZN(_01883_ ) );
BUF_X4 _19723_ ( .A(_04731_ ), .Z(_05037_ ) );
NAND4_X1 _19724_ ( .A1(_10632_ ), .A2(_05027_ ), .A3(_05037_ ), .A4(_05005_ ), .ZN(_05038_ ) );
OAI21_X1 _19725_ ( .A(\u_lsu.pmem[1478] ), .B1(_02814_ ), .B2(_05019_ ), .ZN(_05039_ ) );
AOI21_X1 _19726_ ( .A(fanout_net_65 ), .B1(_05038_ ), .B2(_05039_ ), .ZN(_01884_ ) );
NAND4_X1 _19727_ ( .A1(_10635_ ), .A2(_05027_ ), .A3(_05037_ ), .A4(_05005_ ), .ZN(_05040_ ) );
OAI21_X1 _19728_ ( .A(\u_lsu.pmem[1477] ), .B1(_02814_ ), .B2(_05019_ ), .ZN(_05041_ ) );
AOI21_X1 _19729_ ( .A(fanout_net_65 ), .B1(_05040_ ), .B2(_05041_ ), .ZN(_01885_ ) );
BUF_X4 _19730_ ( .A(_04685_ ), .Z(_05042_ ) );
NAND4_X1 _19731_ ( .A1(_10641_ ), .A2(_05027_ ), .A3(_05037_ ), .A4(_05042_ ), .ZN(_05043_ ) );
OAI21_X1 _19732_ ( .A(\u_lsu.pmem[1476] ), .B1(_02814_ ), .B2(_05019_ ), .ZN(_05044_ ) );
AOI21_X1 _19733_ ( .A(fanout_net_65 ), .B1(_05043_ ), .B2(_05044_ ), .ZN(_01886_ ) );
NAND4_X1 _19734_ ( .A1(_10645_ ), .A2(_05027_ ), .A3(_05037_ ), .A4(_05042_ ), .ZN(_05045_ ) );
BUF_X8 _19735_ ( .A(_09450_ ), .Z(_05046_ ) );
BUF_X4 _19736_ ( .A(_05046_ ), .Z(_05047_ ) );
OAI21_X1 _19737_ ( .A(\u_lsu.pmem[1475] ), .B1(_02814_ ), .B2(_05047_ ), .ZN(_05048_ ) );
AOI21_X1 _19738_ ( .A(fanout_net_65 ), .B1(_05045_ ), .B2(_05048_ ), .ZN(_01887_ ) );
NAND2_X1 _19739_ ( .A1(_04941_ ), .A2(\u_lsu.pmem[4099] ), .ZN(_05049_ ) );
NAND4_X1 _19740_ ( .A1(_04669_ ), .A2(_09519_ ), .A3(_10589_ ), .A4(_02485_ ), .ZN(_05050_ ) );
AOI21_X1 _19741_ ( .A(fanout_net_65 ), .B1(_05049_ ), .B2(_05050_ ), .ZN(_01888_ ) );
NAND4_X1 _19742_ ( .A1(_10649_ ), .A2(_05027_ ), .A3(_05037_ ), .A4(_05042_ ), .ZN(_05051_ ) );
OAI21_X1 _19743_ ( .A(\u_lsu.pmem[1474] ), .B1(_02814_ ), .B2(_05047_ ), .ZN(_05052_ ) );
AOI21_X1 _19744_ ( .A(fanout_net_65 ), .B1(_05051_ ), .B2(_05052_ ), .ZN(_01889_ ) );
NAND4_X1 _19745_ ( .A1(_10652_ ), .A2(_05030_ ), .A3(_05037_ ), .A4(_05042_ ), .ZN(_05053_ ) );
OAI21_X1 _19746_ ( .A(\u_lsu.pmem[1473] ), .B1(_02814_ ), .B2(_05047_ ), .ZN(_05054_ ) );
AOI21_X1 _19747_ ( .A(fanout_net_65 ), .B1(_05053_ ), .B2(_05054_ ), .ZN(_01890_ ) );
NAND4_X1 _19748_ ( .A1(_10655_ ), .A2(_05027_ ), .A3(_05037_ ), .A4(_05042_ ), .ZN(_05055_ ) );
OAI21_X1 _19749_ ( .A(\u_lsu.pmem[1472] ), .B1(_02814_ ), .B2(_05047_ ), .ZN(_05056_ ) );
AOI21_X1 _19750_ ( .A(fanout_net_65 ), .B1(_05055_ ), .B2(_05056_ ), .ZN(_01891_ ) );
NAND4_X1 _19751_ ( .A1(_10658_ ), .A2(_05027_ ), .A3(_05037_ ), .A4(_05042_ ), .ZN(_05057_ ) );
OAI21_X1 _19752_ ( .A(\u_lsu.pmem[1447] ), .B1(_02839_ ), .B2(_05047_ ), .ZN(_05058_ ) );
AOI21_X1 _19753_ ( .A(fanout_net_65 ), .B1(_05057_ ), .B2(_05058_ ), .ZN(_01892_ ) );
NAND4_X1 _19754_ ( .A1(_10665_ ), .A2(_05030_ ), .A3(_05037_ ), .A4(_05042_ ), .ZN(_05059_ ) );
OAI21_X1 _19755_ ( .A(\u_lsu.pmem[1446] ), .B1(_02839_ ), .B2(_05047_ ), .ZN(_05060_ ) );
AOI21_X1 _19756_ ( .A(fanout_net_65 ), .B1(_05059_ ), .B2(_05060_ ), .ZN(_01893_ ) );
NAND4_X1 _19757_ ( .A1(_10668_ ), .A2(_05027_ ), .A3(_05037_ ), .A4(_05042_ ), .ZN(_05061_ ) );
OAI21_X1 _19758_ ( .A(\u_lsu.pmem[1445] ), .B1(_02839_ ), .B2(_05047_ ), .ZN(_05062_ ) );
AOI21_X1 _19759_ ( .A(fanout_net_65 ), .B1(_05061_ ), .B2(_05062_ ), .ZN(_01894_ ) );
BUF_X4 _19760_ ( .A(_04731_ ), .Z(_05063_ ) );
NAND4_X1 _19761_ ( .A1(_10671_ ), .A2(_05030_ ), .A3(_05063_ ), .A4(_05042_ ), .ZN(_05064_ ) );
OAI21_X1 _19762_ ( .A(\u_lsu.pmem[1444] ), .B1(_02839_ ), .B2(_05047_ ), .ZN(_05065_ ) );
AOI21_X1 _19763_ ( .A(fanout_net_65 ), .B1(_05064_ ), .B2(_05065_ ), .ZN(_01895_ ) );
NAND4_X1 _19764_ ( .A1(_10674_ ), .A2(_05030_ ), .A3(_05063_ ), .A4(_05042_ ), .ZN(_05066_ ) );
OAI21_X1 _19765_ ( .A(\u_lsu.pmem[1443] ), .B1(_02839_ ), .B2(_05047_ ), .ZN(_05067_ ) );
AOI21_X1 _19766_ ( .A(fanout_net_65 ), .B1(_05066_ ), .B2(_05067_ ), .ZN(_01896_ ) );
BUF_X4 _19767_ ( .A(_04685_ ), .Z(_05068_ ) );
NAND4_X1 _19768_ ( .A1(_10679_ ), .A2(_05030_ ), .A3(_05063_ ), .A4(_05068_ ), .ZN(_05069_ ) );
OAI21_X1 _19769_ ( .A(\u_lsu.pmem[1442] ), .B1(_02839_ ), .B2(_05047_ ), .ZN(_05070_ ) );
AOI21_X1 _19770_ ( .A(fanout_net_65 ), .B1(_05069_ ), .B2(_05070_ ), .ZN(_01897_ ) );
NAND4_X1 _19771_ ( .A1(_10682_ ), .A2(_05030_ ), .A3(_05063_ ), .A4(_05068_ ), .ZN(_05071_ ) );
BUF_X4 _19772_ ( .A(_05046_ ), .Z(_05072_ ) );
OAI21_X1 _19773_ ( .A(\u_lsu.pmem[1441] ), .B1(_02839_ ), .B2(_05072_ ), .ZN(_05073_ ) );
AOI21_X1 _19774_ ( .A(fanout_net_65 ), .B1(_05071_ ), .B2(_05073_ ), .ZN(_01898_ ) );
NAND3_X1 _19775_ ( .A1(_11021_ ), .A2(_10064_ ), .A3(_11212_ ), .ZN(_05074_ ) );
NAND2_X1 _19776_ ( .A1(_04941_ ), .A2(\u_lsu.pmem[4098] ), .ZN(_05075_ ) );
AOI21_X1 _19777_ ( .A(fanout_net_65 ), .B1(_05074_ ), .B2(_05075_ ), .ZN(_01899_ ) );
NAND4_X1 _19778_ ( .A1(_04987_ ), .A2(_04964_ ), .A3(_03753_ ), .A4(_10661_ ), .ZN(_05076_ ) );
OAI21_X1 _19779_ ( .A(\u_lsu.pmem[1440] ), .B1(_02839_ ), .B2(_05072_ ), .ZN(_05077_ ) );
AOI21_X1 _19780_ ( .A(fanout_net_65 ), .B1(_05076_ ), .B2(_05077_ ), .ZN(_01900_ ) );
OAI21_X1 _19781_ ( .A(\u_lsu.pmem[1415] ), .B1(_02860_ ), .B2(_04593_ ), .ZN(_05078_ ) );
NAND4_X1 _19782_ ( .A1(_10694_ ), .A2(_03478_ ), .A3(_04862_ ), .A4(_04595_ ), .ZN(_05079_ ) );
AOI21_X1 _19783_ ( .A(fanout_net_65 ), .B1(_05078_ ), .B2(_05079_ ), .ZN(_01901_ ) );
OAI21_X1 _19784_ ( .A(\u_lsu.pmem[1414] ), .B1(_02860_ ), .B2(_04593_ ), .ZN(_05080_ ) );
NAND4_X1 _19785_ ( .A1(_10694_ ), .A2(_09575_ ), .A3(_04862_ ), .A4(_04595_ ), .ZN(_05081_ ) );
AOI21_X1 _19786_ ( .A(fanout_net_65 ), .B1(_05080_ ), .B2(_05081_ ), .ZN(_01902_ ) );
OAI21_X1 _19787_ ( .A(\u_lsu.pmem[1413] ), .B1(_02859_ ), .B2(_04593_ ), .ZN(_05082_ ) );
NAND4_X1 _19788_ ( .A1(_10694_ ), .A2(_09582_ ), .A3(_04862_ ), .A4(_04595_ ), .ZN(_05083_ ) );
AOI21_X1 _19789_ ( .A(fanout_net_65 ), .B1(_05082_ ), .B2(_05083_ ), .ZN(_01903_ ) );
BUF_X4 _19790_ ( .A(_10720_ ), .Z(_05084_ ) );
OAI21_X1 _19791_ ( .A(\u_lsu.pmem[1412] ), .B1(_02859_ ), .B2(_05084_ ), .ZN(_05085_ ) );
BUF_X4 _19792_ ( .A(_09522_ ), .Z(_05086_ ) );
NAND4_X1 _19793_ ( .A1(_10694_ ), .A2(_08605_ ), .A3(_04862_ ), .A4(_05086_ ), .ZN(_05087_ ) );
AOI21_X1 _19794_ ( .A(fanout_net_65 ), .B1(_05085_ ), .B2(_05087_ ), .ZN(_01904_ ) );
OAI21_X1 _19795_ ( .A(\u_lsu.pmem[1411] ), .B1(_02859_ ), .B2(_05084_ ), .ZN(_05088_ ) );
NAND4_X1 _19796_ ( .A1(_10694_ ), .A2(_09519_ ), .A3(_04862_ ), .A4(_05086_ ), .ZN(_05089_ ) );
AOI21_X1 _19797_ ( .A(fanout_net_65 ), .B1(_05088_ ), .B2(_05089_ ), .ZN(_01905_ ) );
OAI21_X1 _19798_ ( .A(\u_lsu.pmem[1410] ), .B1(_02859_ ), .B2(_05084_ ), .ZN(_05090_ ) );
NAND4_X1 _19799_ ( .A1(_09537_ ), .A2(_10126_ ), .A3(_04862_ ), .A4(_05086_ ), .ZN(_05091_ ) );
AOI21_X1 _19800_ ( .A(fanout_net_65 ), .B1(_05090_ ), .B2(_05091_ ), .ZN(_01906_ ) );
OAI21_X1 _19801_ ( .A(\u_lsu.pmem[1409] ), .B1(_02859_ ), .B2(_05084_ ), .ZN(_05092_ ) );
BUF_X4 _19802_ ( .A(_09455_ ), .Z(_05093_ ) );
NAND4_X1 _19803_ ( .A1(_10694_ ), .A2(_09543_ ), .A3(_05093_ ), .A4(_05086_ ), .ZN(_05094_ ) );
AOI21_X1 _19804_ ( .A(fanout_net_65 ), .B1(_05092_ ), .B2(_05094_ ), .ZN(_01907_ ) );
OAI21_X1 _19805_ ( .A(\u_lsu.pmem[1408] ), .B1(_02859_ ), .B2(_05084_ ), .ZN(_05095_ ) );
NAND4_X1 _19806_ ( .A1(_10694_ ), .A2(_09547_ ), .A3(_05093_ ), .A4(_05086_ ), .ZN(_05096_ ) );
AOI21_X1 _19807_ ( .A(fanout_net_65 ), .B1(_05095_ ), .B2(_05096_ ), .ZN(_01908_ ) );
NAND3_X1 _19808_ ( .A1(_05008_ ), .A2(_11138_ ), .A3(_02884_ ), .ZN(_05097_ ) );
OAI21_X1 _19809_ ( .A(\u_lsu.pmem[1383] ), .B1(_04997_ ), .B2(_02888_ ), .ZN(_05098_ ) );
AOI21_X1 _19810_ ( .A(fanout_net_65 ), .B1(_05097_ ), .B2(_05098_ ), .ZN(_01909_ ) );
NAND2_X1 _19811_ ( .A1(_04941_ ), .A2(\u_lsu.pmem[4097] ), .ZN(_05099_ ) );
NAND4_X1 _19812_ ( .A1(_04669_ ), .A2(_09543_ ), .A3(_10589_ ), .A4(_02485_ ), .ZN(_05100_ ) );
AOI21_X1 _19813_ ( .A(fanout_net_65 ), .B1(_05099_ ), .B2(_05100_ ), .ZN(_01910_ ) );
NAND4_X1 _19814_ ( .A1(_04987_ ), .A2(_09925_ ), .A3(_05063_ ), .A4(_03786_ ), .ZN(_05101_ ) );
OAI21_X1 _19815_ ( .A(\u_lsu.pmem[1382] ), .B1(_04997_ ), .B2(_02888_ ), .ZN(_05102_ ) );
AOI21_X1 _19816_ ( .A(fanout_net_66 ), .B1(_05101_ ), .B2(_05102_ ), .ZN(_01911_ ) );
NAND4_X1 _19817_ ( .A1(_04987_ ), .A2(_09928_ ), .A3(_05063_ ), .A4(_03786_ ), .ZN(_05103_ ) );
OAI21_X1 _19818_ ( .A(\u_lsu.pmem[1381] ), .B1(_04997_ ), .B2(_02888_ ), .ZN(_05104_ ) );
AOI21_X1 _19819_ ( .A(fanout_net_66 ), .B1(_05103_ ), .B2(_05104_ ), .ZN(_01912_ ) );
NAND4_X1 _19820_ ( .A1(_04987_ ), .A2(_09931_ ), .A3(_05063_ ), .A4(_03786_ ), .ZN(_05105_ ) );
BUF_X4 _19821_ ( .A(_04571_ ), .Z(_05106_ ) );
OAI21_X1 _19822_ ( .A(\u_lsu.pmem[1380] ), .B1(_05106_ ), .B2(_02885_ ), .ZN(_05107_ ) );
AOI21_X1 _19823_ ( .A(fanout_net_66 ), .B1(_05105_ ), .B2(_05107_ ), .ZN(_01913_ ) );
NAND4_X1 _19824_ ( .A1(_04987_ ), .A2(_03091_ ), .A3(_05063_ ), .A4(_03786_ ), .ZN(_05108_ ) );
OAI21_X1 _19825_ ( .A(\u_lsu.pmem[1379] ), .B1(_05106_ ), .B2(_02885_ ), .ZN(_05109_ ) );
AOI21_X1 _19826_ ( .A(fanout_net_66 ), .B1(_05108_ ), .B2(_05109_ ), .ZN(_01914_ ) );
NAND4_X1 _19827_ ( .A1(_04987_ ), .A2(_09938_ ), .A3(_05063_ ), .A4(_03786_ ), .ZN(_05110_ ) );
OAI21_X1 _19828_ ( .A(\u_lsu.pmem[1378] ), .B1(_05106_ ), .B2(_02885_ ), .ZN(_05111_ ) );
AOI21_X1 _19829_ ( .A(fanout_net_66 ), .B1(_05110_ ), .B2(_05111_ ), .ZN(_01915_ ) );
NAND4_X1 _19830_ ( .A1(_04987_ ), .A2(_03143_ ), .A3(_05063_ ), .A4(_03786_ ), .ZN(_05112_ ) );
OAI21_X1 _19831_ ( .A(\u_lsu.pmem[1377] ), .B1(_05106_ ), .B2(_02885_ ), .ZN(_05113_ ) );
AOI21_X1 _19832_ ( .A(fanout_net_66 ), .B1(_05112_ ), .B2(_05113_ ), .ZN(_01916_ ) );
BUF_X4 _19833_ ( .A(_10036_ ), .Z(_05114_ ) );
BUF_X4 _19834_ ( .A(_04731_ ), .Z(_05115_ ) );
NAND4_X1 _19835_ ( .A1(_05114_ ), .A2(_09944_ ), .A3(_05115_ ), .A4(_10723_ ), .ZN(_05116_ ) );
OAI21_X1 _19836_ ( .A(\u_lsu.pmem[1376] ), .B1(_05106_ ), .B2(_02885_ ), .ZN(_05117_ ) );
AOI21_X1 _19837_ ( .A(fanout_net_66 ), .B1(_05116_ ), .B2(_05117_ ), .ZN(_01917_ ) );
NAND3_X1 _19838_ ( .A1(_05008_ ), .A2(_11138_ ), .A3(_02908_ ), .ZN(_05118_ ) );
OAI21_X1 _19839_ ( .A(\u_lsu.pmem[1351] ), .B1(_05106_ ), .B2(_02910_ ), .ZN(_05119_ ) );
AOI21_X1 _19840_ ( .A(fanout_net_66 ), .B1(_05118_ ), .B2(_05119_ ), .ZN(_01918_ ) );
NAND4_X1 _19841_ ( .A1(_05114_ ), .A2(_09925_ ), .A3(_05115_ ), .A4(_03804_ ), .ZN(_05120_ ) );
OAI21_X1 _19842_ ( .A(\u_lsu.pmem[1350] ), .B1(_05106_ ), .B2(_02910_ ), .ZN(_05121_ ) );
AOI21_X1 _19843_ ( .A(fanout_net_66 ), .B1(_05120_ ), .B2(_05121_ ), .ZN(_01919_ ) );
NAND4_X1 _19844_ ( .A1(_05114_ ), .A2(_09928_ ), .A3(_05115_ ), .A4(_03804_ ), .ZN(_05122_ ) );
OAI21_X1 _19845_ ( .A(\u_lsu.pmem[1349] ), .B1(_05106_ ), .B2(_02909_ ), .ZN(_05123_ ) );
AOI21_X1 _19846_ ( .A(fanout_net_66 ), .B1(_05122_ ), .B2(_05123_ ), .ZN(_01920_ ) );
NAND2_X1 _19847_ ( .A1(_04941_ ), .A2(\u_lsu.pmem[4096] ), .ZN(_05124_ ) );
NAND4_X1 _19848_ ( .A1(_04669_ ), .A2(_09547_ ), .A3(_10046_ ), .A4(_02485_ ), .ZN(_05125_ ) );
AOI21_X1 _19849_ ( .A(fanout_net_66 ), .B1(_05124_ ), .B2(_05125_ ), .ZN(_01921_ ) );
NAND4_X1 _19850_ ( .A1(_05114_ ), .A2(_09931_ ), .A3(_05115_ ), .A4(_03804_ ), .ZN(_05126_ ) );
OAI21_X1 _19851_ ( .A(\u_lsu.pmem[1348] ), .B1(_05106_ ), .B2(_02909_ ), .ZN(_05127_ ) );
AOI21_X1 _19852_ ( .A(fanout_net_66 ), .B1(_05126_ ), .B2(_05127_ ), .ZN(_01922_ ) );
NAND4_X1 _19853_ ( .A1(_05114_ ), .A2(_03091_ ), .A3(_05115_ ), .A4(_03804_ ), .ZN(_05128_ ) );
OAI21_X1 _19854_ ( .A(\u_lsu.pmem[1347] ), .B1(_05106_ ), .B2(_02909_ ), .ZN(_05129_ ) );
AOI21_X1 _19855_ ( .A(fanout_net_66 ), .B1(_05128_ ), .B2(_05129_ ), .ZN(_01923_ ) );
NAND4_X1 _19856_ ( .A1(_05114_ ), .A2(_09938_ ), .A3(_05115_ ), .A4(_03804_ ), .ZN(_05130_ ) );
BUF_X4 _19857_ ( .A(_09472_ ), .Z(_05131_ ) );
OAI21_X1 _19858_ ( .A(\u_lsu.pmem[1346] ), .B1(_05131_ ), .B2(_02909_ ), .ZN(_05132_ ) );
AOI21_X1 _19859_ ( .A(fanout_net_66 ), .B1(_05130_ ), .B2(_05132_ ), .ZN(_01924_ ) );
NAND4_X1 _19860_ ( .A1(_05114_ ), .A2(_03143_ ), .A3(_05115_ ), .A4(_10750_ ), .ZN(_05133_ ) );
OAI21_X1 _19861_ ( .A(\u_lsu.pmem[1345] ), .B1(_05131_ ), .B2(_02909_ ), .ZN(_05134_ ) );
AOI21_X1 _19862_ ( .A(fanout_net_66 ), .B1(_05133_ ), .B2(_05134_ ), .ZN(_01925_ ) );
NAND4_X1 _19863_ ( .A1(_05114_ ), .A2(_09944_ ), .A3(_05115_ ), .A4(_10750_ ), .ZN(_05135_ ) );
OAI21_X1 _19864_ ( .A(\u_lsu.pmem[1344] ), .B1(_05131_ ), .B2(_02909_ ), .ZN(_05136_ ) );
AOI21_X1 _19865_ ( .A(fanout_net_66 ), .B1(_05135_ ), .B2(_05136_ ), .ZN(_01926_ ) );
NAND4_X1 _19866_ ( .A1(_09670_ ), .A2(_05030_ ), .A3(_05115_ ), .A4(_05068_ ), .ZN(_05137_ ) );
OAI21_X1 _19867_ ( .A(\u_lsu.pmem[1319] ), .B1(_02932_ ), .B2(_05072_ ), .ZN(_05138_ ) );
AOI21_X1 _19868_ ( .A(fanout_net_66 ), .B1(_05137_ ), .B2(_05138_ ), .ZN(_01927_ ) );
NAND4_X1 _19869_ ( .A1(_09681_ ), .A2(_05030_ ), .A3(_05115_ ), .A4(_05068_ ), .ZN(_05139_ ) );
OAI21_X1 _19870_ ( .A(\u_lsu.pmem[1318] ), .B1(_02932_ ), .B2(_05072_ ), .ZN(_05140_ ) );
AOI21_X1 _19871_ ( .A(fanout_net_66 ), .B1(_05139_ ), .B2(_05140_ ), .ZN(_01928_ ) );
BUF_X4 _19872_ ( .A(_04731_ ), .Z(_05141_ ) );
NAND4_X1 _19873_ ( .A1(_09685_ ), .A2(_05030_ ), .A3(_05141_ ), .A4(_05068_ ), .ZN(_05142_ ) );
OAI21_X1 _19874_ ( .A(\u_lsu.pmem[1317] ), .B1(_02932_ ), .B2(_05072_ ), .ZN(_05143_ ) );
AOI21_X1 _19875_ ( .A(fanout_net_66 ), .B1(_05142_ ), .B2(_05143_ ), .ZN(_01929_ ) );
AND3_X1 _19876_ ( .A1(_09149_ ), .A2(_04008_ ), .A3(_02931_ ), .ZN(_05144_ ) );
AOI21_X1 _19877_ ( .A(\u_lsu.pmem[1316] ), .B1(_09676_ ), .B2(_02931_ ), .ZN(_05145_ ) );
NOR3_X1 _19878_ ( .A1(_05144_ ), .A2(_05145_ ), .A3(fanout_net_66 ), .ZN(_01930_ ) );
OAI21_X1 _19879_ ( .A(\u_lsu.pmem[1315] ), .B1(_02933_ ), .B2(_05084_ ), .ZN(_05146_ ) );
NAND3_X1 _19880_ ( .A1(_04470_ ), .A2(_02931_ ), .A3(_09449_ ), .ZN(_05147_ ) );
AOI21_X1 _19881_ ( .A(fanout_net_66 ), .B1(_05146_ ), .B2(_05147_ ), .ZN(_01931_ ) );
AND2_X1 _19882_ ( .A1(_10057_ ), .A2(_10012_ ), .ZN(_05148_ ) );
OAI21_X1 _19883_ ( .A(_09109_ ), .B1(_05148_ ), .B2(\u_lsu.pmem[4071] ), .ZN(_05149_ ) );
AOI21_X1 _19884_ ( .A(_05149_ ), .B1(_09568_ ), .B2(_05148_ ), .ZN(_01932_ ) );
OAI21_X1 _19885_ ( .A(\u_lsu.pmem[1314] ), .B1(_02933_ ), .B2(_05084_ ), .ZN(_05150_ ) );
NAND3_X1 _19886_ ( .A1(_04470_ ), .A2(_02931_ ), .A3(_10492_ ), .ZN(_05151_ ) );
AOI21_X1 _19887_ ( .A(fanout_net_66 ), .B1(_05150_ ), .B2(_05151_ ), .ZN(_01933_ ) );
OAI21_X1 _19888_ ( .A(\u_lsu.pmem[1313] ), .B1(_02933_ ), .B2(_05084_ ), .ZN(_05152_ ) );
NAND3_X1 _19889_ ( .A1(_04470_ ), .A2(_02931_ ), .A3(_09698_ ), .ZN(_05153_ ) );
AOI21_X1 _19890_ ( .A(fanout_net_66 ), .B1(_05152_ ), .B2(_05153_ ), .ZN(_01934_ ) );
BUF_X4 _19891_ ( .A(_10063_ ), .Z(_05154_ ) );
NAND4_X1 _19892_ ( .A1(_09703_ ), .A2(_05154_ ), .A3(_05141_ ), .A4(_05068_ ), .ZN(_05155_ ) );
OAI21_X1 _19893_ ( .A(\u_lsu.pmem[1312] ), .B1(_02932_ ), .B2(_05072_ ), .ZN(_05156_ ) );
AOI21_X1 _19894_ ( .A(fanout_net_66 ), .B1(_05155_ ), .B2(_05156_ ), .ZN(_01935_ ) );
BUF_X4 _19895_ ( .A(_10287_ ), .Z(_05157_ ) );
NAND4_X1 _19896_ ( .A1(_09708_ ), .A2(_05157_ ), .A3(_05141_ ), .A4(_05068_ ), .ZN(_05158_ ) );
OAI21_X1 _19897_ ( .A(\u_lsu.pmem[1287] ), .B1(_02957_ ), .B2(_05072_ ), .ZN(_05159_ ) );
AOI21_X1 _19898_ ( .A(fanout_net_66 ), .B1(_05158_ ), .B2(_05159_ ), .ZN(_01936_ ) );
NAND4_X1 _19899_ ( .A1(_09715_ ), .A2(_05157_ ), .A3(_05141_ ), .A4(_05068_ ), .ZN(_05160_ ) );
OAI21_X1 _19900_ ( .A(\u_lsu.pmem[1286] ), .B1(_02957_ ), .B2(_05072_ ), .ZN(_05161_ ) );
AOI21_X1 _19901_ ( .A(fanout_net_66 ), .B1(_05160_ ), .B2(_05161_ ), .ZN(_01937_ ) );
NAND4_X1 _19902_ ( .A1(_09718_ ), .A2(_05157_ ), .A3(_05141_ ), .A4(_05068_ ), .ZN(_05162_ ) );
OAI21_X1 _19903_ ( .A(\u_lsu.pmem[1285] ), .B1(_02957_ ), .B2(_05072_ ), .ZN(_05163_ ) );
AOI21_X1 _19904_ ( .A(fanout_net_66 ), .B1(_05162_ ), .B2(_05163_ ), .ZN(_01938_ ) );
NAND4_X1 _19905_ ( .A1(_09721_ ), .A2(_05157_ ), .A3(_05141_ ), .A4(_05068_ ), .ZN(_05164_ ) );
OAI21_X1 _19906_ ( .A(\u_lsu.pmem[1284] ), .B1(_02957_ ), .B2(_05072_ ), .ZN(_05165_ ) );
AOI21_X1 _19907_ ( .A(fanout_net_66 ), .B1(_05164_ ), .B2(_05165_ ), .ZN(_01939_ ) );
BUF_X8 _19908_ ( .A(_09442_ ), .Z(_05166_ ) );
BUF_X4 _19909_ ( .A(_05166_ ), .Z(_05167_ ) );
NAND4_X1 _19910_ ( .A1(_09725_ ), .A2(_05157_ ), .A3(_05141_ ), .A4(_05167_ ), .ZN(_05168_ ) );
BUF_X4 _19911_ ( .A(_05046_ ), .Z(_05169_ ) );
OAI21_X1 _19912_ ( .A(\u_lsu.pmem[1283] ), .B1(_02957_ ), .B2(_05169_ ), .ZN(_05170_ ) );
AOI21_X1 _19913_ ( .A(fanout_net_66 ), .B1(_05168_ ), .B2(_05170_ ), .ZN(_01940_ ) );
NAND4_X1 _19914_ ( .A1(_05114_ ), .A2(_09474_ ), .A3(_05141_ ), .A4(_10797_ ), .ZN(_05171_ ) );
OAI21_X1 _19915_ ( .A(\u_lsu.pmem[1282] ), .B1(_02957_ ), .B2(_05169_ ), .ZN(_05172_ ) );
AOI21_X1 _19916_ ( .A(fanout_net_66 ), .B1(_05171_ ), .B2(_05172_ ), .ZN(_01941_ ) );
NAND4_X1 _19917_ ( .A1(_09733_ ), .A2(_05154_ ), .A3(_05141_ ), .A4(_05167_ ), .ZN(_05173_ ) );
OAI21_X1 _19918_ ( .A(\u_lsu.pmem[1281] ), .B1(_02957_ ), .B2(_05169_ ), .ZN(_05174_ ) );
AOI21_X1 _19919_ ( .A(fanout_net_67 ), .B1(_05173_ ), .B2(_05174_ ), .ZN(_01942_ ) );
NAND4_X1 _19920_ ( .A1(_10062_ ), .A2(_05154_ ), .A3(_04658_ ), .A4(_05167_ ), .ZN(_05175_ ) );
OAI21_X1 _19921_ ( .A(\u_lsu.pmem[4070] ), .B1(_10069_ ), .B2(_04671_ ), .ZN(_05176_ ) );
AOI21_X1 _19922_ ( .A(fanout_net_67 ), .B1(_05175_ ), .B2(_05176_ ), .ZN(_01943_ ) );
NAND4_X1 _19923_ ( .A1(_09736_ ), .A2(_05157_ ), .A3(_05141_ ), .A4(_05167_ ), .ZN(_05177_ ) );
OAI21_X1 _19924_ ( .A(\u_lsu.pmem[1280] ), .B1(_02957_ ), .B2(_05169_ ), .ZN(_05178_ ) );
AOI21_X1 _19925_ ( .A(fanout_net_67 ), .B1(_05177_ ), .B2(_05178_ ), .ZN(_01944_ ) );
NAND4_X1 _19926_ ( .A1(_05114_ ), .A2(_04964_ ), .A3(_04928_ ), .A4(_10819_ ), .ZN(_05179_ ) );
OAI21_X1 _19927_ ( .A(\u_lsu.pmem[1255] ), .B1(_02982_ ), .B2(_05169_ ), .ZN(_05180_ ) );
AOI21_X1 _19928_ ( .A(fanout_net_67 ), .B1(_05179_ ), .B2(_05180_ ), .ZN(_01945_ ) );
BUF_X8 _19929_ ( .A(_09455_ ), .Z(_05181_ ) );
BUF_X4 _19930_ ( .A(_05181_ ), .Z(_05182_ ) );
NAND4_X1 _19931_ ( .A1(_09756_ ), .A2(_05157_ ), .A3(_05182_ ), .A4(_05167_ ), .ZN(_05183_ ) );
OAI21_X1 _19932_ ( .A(\u_lsu.pmem[1254] ), .B1(_02982_ ), .B2(_05169_ ), .ZN(_05184_ ) );
AOI21_X1 _19933_ ( .A(fanout_net_67 ), .B1(_05183_ ), .B2(_05184_ ), .ZN(_01946_ ) );
NAND4_X1 _19934_ ( .A1(_09763_ ), .A2(_05154_ ), .A3(_05182_ ), .A4(_05167_ ), .ZN(_05185_ ) );
OAI21_X1 _19935_ ( .A(\u_lsu.pmem[1253] ), .B1(_02982_ ), .B2(_05169_ ), .ZN(_05186_ ) );
AOI21_X1 _19936_ ( .A(fanout_net_67 ), .B1(_05185_ ), .B2(_05186_ ), .ZN(_01947_ ) );
NAND4_X1 _19937_ ( .A1(_09770_ ), .A2(_05157_ ), .A3(_05182_ ), .A4(_05167_ ), .ZN(_05187_ ) );
OAI21_X1 _19938_ ( .A(\u_lsu.pmem[1252] ), .B1(_02982_ ), .B2(_05169_ ), .ZN(_05188_ ) );
AOI21_X1 _19939_ ( .A(fanout_net_67 ), .B1(_05187_ ), .B2(_05188_ ), .ZN(_01948_ ) );
NAND4_X1 _19940_ ( .A1(_09775_ ), .A2(_05154_ ), .A3(_05182_ ), .A4(_05167_ ), .ZN(_05189_ ) );
OAI21_X1 _19941_ ( .A(\u_lsu.pmem[1251] ), .B1(_02982_ ), .B2(_05169_ ), .ZN(_05190_ ) );
AOI21_X1 _19942_ ( .A(fanout_net_67 ), .B1(_05189_ ), .B2(_05190_ ), .ZN(_01949_ ) );
NAND4_X1 _19943_ ( .A1(_09780_ ), .A2(_05154_ ), .A3(_05182_ ), .A4(_05167_ ), .ZN(_05191_ ) );
OAI21_X1 _19944_ ( .A(\u_lsu.pmem[1250] ), .B1(_02982_ ), .B2(_05169_ ), .ZN(_05192_ ) );
AOI21_X1 _19945_ ( .A(fanout_net_67 ), .B1(_05191_ ), .B2(_05192_ ), .ZN(_01950_ ) );
NAND4_X1 _19946_ ( .A1(_09787_ ), .A2(_05154_ ), .A3(_05182_ ), .A4(_05167_ ), .ZN(_05193_ ) );
BUF_X4 _19947_ ( .A(_05046_ ), .Z(_05194_ ) );
OAI21_X1 _19948_ ( .A(\u_lsu.pmem[1249] ), .B1(_02982_ ), .B2(_05194_ ), .ZN(_05195_ ) );
AOI21_X1 _19949_ ( .A(fanout_net_67 ), .B1(_05193_ ), .B2(_05195_ ), .ZN(_01951_ ) );
BUF_X4 _19950_ ( .A(_05166_ ), .Z(_05196_ ) );
NAND4_X1 _19951_ ( .A1(_09791_ ), .A2(_05154_ ), .A3(_05182_ ), .A4(_05196_ ), .ZN(_05197_ ) );
OAI21_X1 _19952_ ( .A(\u_lsu.pmem[1248] ), .B1(_02982_ ), .B2(_05194_ ), .ZN(_05198_ ) );
AOI21_X1 _19953_ ( .A(fanout_net_67 ), .B1(_05197_ ), .B2(_05198_ ), .ZN(_01952_ ) );
BUF_X4 _19954_ ( .A(_10036_ ), .Z(_05199_ ) );
NAND4_X1 _19955_ ( .A1(_05199_ ), .A2(_09674_ ), .A3(_04928_ ), .A4(_10847_ ), .ZN(_05200_ ) );
OAI21_X1 _19956_ ( .A(\u_lsu.pmem[1223] ), .B1(_03005_ ), .B2(_05194_ ), .ZN(_05201_ ) );
AOI21_X1 _19957_ ( .A(fanout_net_67 ), .B1(_05200_ ), .B2(_05201_ ), .ZN(_01953_ ) );
NAND4_X1 _19958_ ( .A1(_10075_ ), .A2(_05154_ ), .A3(_04658_ ), .A4(_05196_ ), .ZN(_05202_ ) );
OAI21_X1 _19959_ ( .A(\u_lsu.pmem[4069] ), .B1(_10069_ ), .B2(_04671_ ), .ZN(_05203_ ) );
AOI21_X1 _19960_ ( .A(fanout_net_67 ), .B1(_05202_ ), .B2(_05203_ ), .ZN(_01954_ ) );
NAND4_X1 _19961_ ( .A1(_09804_ ), .A2(_02486_ ), .A3(_10585_ ), .A4(_05196_ ), .ZN(_05204_ ) );
OAI21_X1 _19962_ ( .A(\u_lsu.pmem[1222] ), .B1(_03005_ ), .B2(_05194_ ), .ZN(_05205_ ) );
AOI21_X1 _19963_ ( .A(fanout_net_67 ), .B1(_05204_ ), .B2(_05205_ ), .ZN(_01955_ ) );
NAND4_X1 _19964_ ( .A1(_09811_ ), .A2(_05157_ ), .A3(_05182_ ), .A4(_05196_ ), .ZN(_05206_ ) );
OAI21_X1 _19965_ ( .A(\u_lsu.pmem[1221] ), .B1(_03005_ ), .B2(_05194_ ), .ZN(_05207_ ) );
AOI21_X1 _19966_ ( .A(fanout_net_67 ), .B1(_05206_ ), .B2(_05207_ ), .ZN(_01956_ ) );
NAND4_X1 _19967_ ( .A1(_09815_ ), .A2(_05157_ ), .A3(_05182_ ), .A4(_05196_ ), .ZN(_05208_ ) );
OAI21_X1 _19968_ ( .A(\u_lsu.pmem[1220] ), .B1(_03005_ ), .B2(_05194_ ), .ZN(_05209_ ) );
AOI21_X1 _19969_ ( .A(fanout_net_67 ), .B1(_05208_ ), .B2(_05209_ ), .ZN(_01957_ ) );
NAND4_X1 _19970_ ( .A1(_09819_ ), .A2(_10577_ ), .A3(_05182_ ), .A4(_05196_ ), .ZN(_05210_ ) );
OAI21_X1 _19971_ ( .A(\u_lsu.pmem[1219] ), .B1(_03005_ ), .B2(_05194_ ), .ZN(_05211_ ) );
AOI21_X1 _19972_ ( .A(fanout_net_67 ), .B1(_05210_ ), .B2(_05211_ ), .ZN(_01958_ ) );
BUF_X4 _19973_ ( .A(_05181_ ), .Z(_05212_ ) );
NAND4_X1 _19974_ ( .A1(_09827_ ), .A2(_05154_ ), .A3(_05212_ ), .A4(_05196_ ), .ZN(_05213_ ) );
OAI21_X1 _19975_ ( .A(\u_lsu.pmem[1218] ), .B1(_03005_ ), .B2(_05194_ ), .ZN(_05214_ ) );
AOI21_X1 _19976_ ( .A(fanout_net_67 ), .B1(_05213_ ), .B2(_05214_ ), .ZN(_01959_ ) );
BUF_X4 _19977_ ( .A(_10063_ ), .Z(_05215_ ) );
NAND4_X1 _19978_ ( .A1(_09831_ ), .A2(_05215_ ), .A3(_05212_ ), .A4(_05196_ ), .ZN(_05216_ ) );
OAI21_X1 _19979_ ( .A(\u_lsu.pmem[1217] ), .B1(_03005_ ), .B2(_05194_ ), .ZN(_05217_ ) );
AOI21_X1 _19980_ ( .A(fanout_net_67 ), .B1(_05216_ ), .B2(_05217_ ), .ZN(_01960_ ) );
NAND4_X1 _19981_ ( .A1(_09835_ ), .A2(_05215_ ), .A3(_05212_ ), .A4(_05196_ ), .ZN(_05218_ ) );
OAI21_X1 _19982_ ( .A(\u_lsu.pmem[1216] ), .B1(_03005_ ), .B2(_05194_ ), .ZN(_05219_ ) );
AOI21_X1 _19983_ ( .A(fanout_net_67 ), .B1(_05218_ ), .B2(_05219_ ), .ZN(_01961_ ) );
NAND4_X1 _19984_ ( .A1(_09840_ ), .A2(_05215_ ), .A3(_05212_ ), .A4(_05196_ ), .ZN(_05220_ ) );
BUF_X4 _19985_ ( .A(_05046_ ), .Z(_05221_ ) );
OAI21_X1 _19986_ ( .A(\u_lsu.pmem[1191] ), .B1(_03031_ ), .B2(_05221_ ), .ZN(_05222_ ) );
AOI21_X1 _19987_ ( .A(fanout_net_67 ), .B1(_05220_ ), .B2(_05222_ ), .ZN(_01962_ ) );
BUF_X4 _19988_ ( .A(_05166_ ), .Z(_05223_ ) );
NAND4_X1 _19989_ ( .A1(_09849_ ), .A2(_10577_ ), .A3(_05212_ ), .A4(_05223_ ), .ZN(_05224_ ) );
OAI21_X1 _19990_ ( .A(\u_lsu.pmem[1190] ), .B1(_03031_ ), .B2(_05221_ ), .ZN(_05225_ ) );
AOI21_X1 _19991_ ( .A(fanout_net_67 ), .B1(_05224_ ), .B2(_05225_ ), .ZN(_01963_ ) );
NAND4_X1 _19992_ ( .A1(_09853_ ), .A2(_05215_ ), .A3(_05212_ ), .A4(_05223_ ), .ZN(_05226_ ) );
OAI21_X1 _19993_ ( .A(\u_lsu.pmem[1189] ), .B1(_03031_ ), .B2(_05221_ ), .ZN(_05227_ ) );
AOI21_X1 _19994_ ( .A(fanout_net_67 ), .B1(_05226_ ), .B2(_05227_ ), .ZN(_01964_ ) );
NAND4_X1 _19995_ ( .A1(_09721_ ), .A2(_04914_ ), .A3(_05212_ ), .A4(_04097_ ), .ZN(_05228_ ) );
OAI21_X1 _19996_ ( .A(\u_lsu.pmem[4356] ), .B1(_03950_ ), .B2(_09468_ ), .ZN(_05229_ ) );
AOI21_X1 _19997_ ( .A(fanout_net_67 ), .B1(_05228_ ), .B2(_05229_ ), .ZN(_01965_ ) );
NAND4_X1 _19998_ ( .A1(_10079_ ), .A2(_05215_ ), .A3(_04658_ ), .A4(_05223_ ), .ZN(_05230_ ) );
OAI21_X1 _19999_ ( .A(\u_lsu.pmem[4068] ), .B1(_10069_ ), .B2(_04671_ ), .ZN(_05231_ ) );
AOI21_X1 _20000_ ( .A(fanout_net_67 ), .B1(_05230_ ), .B2(_05231_ ), .ZN(_01966_ ) );
NAND4_X1 _20001_ ( .A1(_09858_ ), .A2(_05215_ ), .A3(_05212_ ), .A4(_05223_ ), .ZN(_05232_ ) );
OAI21_X1 _20002_ ( .A(\u_lsu.pmem[1188] ), .B1(_03031_ ), .B2(_05221_ ), .ZN(_05233_ ) );
AOI21_X1 _20003_ ( .A(fanout_net_67 ), .B1(_05232_ ), .B2(_05233_ ), .ZN(_01967_ ) );
NAND4_X1 _20004_ ( .A1(_09861_ ), .A2(_05215_ ), .A3(_05212_ ), .A4(_05223_ ), .ZN(_05234_ ) );
OAI21_X1 _20005_ ( .A(\u_lsu.pmem[1187] ), .B1(_03031_ ), .B2(_05221_ ), .ZN(_05235_ ) );
AOI21_X1 _20006_ ( .A(fanout_net_67 ), .B1(_05234_ ), .B2(_05235_ ), .ZN(_01968_ ) );
NAND4_X1 _20007_ ( .A1(_09864_ ), .A2(_05215_ ), .A3(_05212_ ), .A4(_05223_ ), .ZN(_05236_ ) );
OAI21_X1 _20008_ ( .A(\u_lsu.pmem[1186] ), .B1(_03031_ ), .B2(_05221_ ), .ZN(_05237_ ) );
AOI21_X1 _20009_ ( .A(fanout_net_67 ), .B1(_05236_ ), .B2(_05237_ ), .ZN(_01969_ ) );
BUF_X4 _20010_ ( .A(_05181_ ), .Z(_05238_ ) );
NAND4_X1 _20011_ ( .A1(_09867_ ), .A2(_05215_ ), .A3(_05238_ ), .A4(_05223_ ), .ZN(_05239_ ) );
OAI21_X1 _20012_ ( .A(\u_lsu.pmem[1185] ), .B1(_03031_ ), .B2(_05221_ ), .ZN(_05240_ ) );
AOI21_X1 _20013_ ( .A(fanout_net_67 ), .B1(_05239_ ), .B2(_05240_ ), .ZN(_01970_ ) );
NAND4_X1 _20014_ ( .A1(_09881_ ), .A2(_10577_ ), .A3(_05238_ ), .A4(_05223_ ), .ZN(_05241_ ) );
OAI21_X1 _20015_ ( .A(\u_lsu.pmem[1184] ), .B1(_03031_ ), .B2(_05221_ ), .ZN(_05242_ ) );
AOI21_X1 _20016_ ( .A(fanout_net_67 ), .B1(_05241_ ), .B2(_05242_ ), .ZN(_01971_ ) );
OAI21_X1 _20017_ ( .A(\u_lsu.pmem[1159] ), .B1(_03050_ ), .B2(_05084_ ), .ZN(_05243_ ) );
NAND4_X1 _20018_ ( .A1(_10898_ ), .A2(_08582_ ), .A3(_05093_ ), .A4(_05086_ ), .ZN(_05244_ ) );
AOI21_X1 _20019_ ( .A(fanout_net_68 ), .B1(_05243_ ), .B2(_05244_ ), .ZN(_01972_ ) );
OAI21_X1 _20020_ ( .A(\u_lsu.pmem[1158] ), .B1(_03050_ ), .B2(_05084_ ), .ZN(_05245_ ) );
NAND4_X1 _20021_ ( .A1(_10898_ ), .A2(_09575_ ), .A3(_05093_ ), .A4(_05086_ ), .ZN(_05246_ ) );
AOI21_X1 _20022_ ( .A(fanout_net_68 ), .B1(_05245_ ), .B2(_05246_ ), .ZN(_01973_ ) );
BUF_X4 _20023_ ( .A(_10720_ ), .Z(_05247_ ) );
OAI21_X1 _20024_ ( .A(\u_lsu.pmem[1157] ), .B1(_03049_ ), .B2(_05247_ ), .ZN(_05248_ ) );
NAND4_X1 _20025_ ( .A1(_10898_ ), .A2(_09582_ ), .A3(_05093_ ), .A4(_05086_ ), .ZN(_05249_ ) );
AOI21_X1 _20026_ ( .A(fanout_net_68 ), .B1(_05248_ ), .B2(_05249_ ), .ZN(_01974_ ) );
OAI21_X1 _20027_ ( .A(\u_lsu.pmem[1156] ), .B1(_03049_ ), .B2(_05247_ ), .ZN(_05250_ ) );
NAND4_X1 _20028_ ( .A1(_10898_ ), .A2(_08605_ ), .A3(_05093_ ), .A4(_05086_ ), .ZN(_05251_ ) );
AOI21_X1 _20029_ ( .A(fanout_net_68 ), .B1(_05250_ ), .B2(_05251_ ), .ZN(_01975_ ) );
OAI21_X1 _20030_ ( .A(\u_lsu.pmem[1155] ), .B1(_03049_ ), .B2(_05247_ ), .ZN(_05252_ ) );
NAND4_X1 _20031_ ( .A1(_10898_ ), .A2(_09519_ ), .A3(_05093_ ), .A4(_05086_ ), .ZN(_05253_ ) );
AOI21_X1 _20032_ ( .A(fanout_net_68 ), .B1(_05252_ ), .B2(_05253_ ), .ZN(_01976_ ) );
NAND4_X1 _20033_ ( .A1(_10084_ ), .A2(_05215_ ), .A3(_04658_ ), .A4(_05223_ ), .ZN(_05254_ ) );
OAI21_X1 _20034_ ( .A(\u_lsu.pmem[4067] ), .B1(_10068_ ), .B2(_04671_ ), .ZN(_05255_ ) );
AOI21_X1 _20035_ ( .A(fanout_net_68 ), .B1(_05254_ ), .B2(_05255_ ), .ZN(_01977_ ) );
OAI21_X1 _20036_ ( .A(\u_lsu.pmem[1154] ), .B1(_03049_ ), .B2(_05247_ ), .ZN(_05256_ ) );
BUF_X4 _20037_ ( .A(_09522_ ), .Z(_05257_ ) );
NAND4_X1 _20038_ ( .A1(_09906_ ), .A2(_10126_ ), .A3(_05093_ ), .A4(_05257_ ), .ZN(_05258_ ) );
AOI21_X1 _20039_ ( .A(fanout_net_68 ), .B1(_05256_ ), .B2(_05258_ ), .ZN(_01978_ ) );
OAI21_X1 _20040_ ( .A(\u_lsu.pmem[1153] ), .B1(_03049_ ), .B2(_05247_ ), .ZN(_05259_ ) );
NAND4_X1 _20041_ ( .A1(_10898_ ), .A2(_09543_ ), .A3(_05093_ ), .A4(_05257_ ), .ZN(_05260_ ) );
AOI21_X1 _20042_ ( .A(fanout_net_68 ), .B1(_05259_ ), .B2(_05260_ ), .ZN(_01979_ ) );
OAI21_X1 _20043_ ( .A(\u_lsu.pmem[1152] ), .B1(_03049_ ), .B2(_05247_ ), .ZN(_05261_ ) );
NAND4_X1 _20044_ ( .A1(_10898_ ), .A2(_09547_ ), .A3(_05093_ ), .A4(_05257_ ), .ZN(_05262_ ) );
AOI21_X1 _20045_ ( .A(fanout_net_68 ), .B1(_05261_ ), .B2(_05262_ ), .ZN(_01980_ ) );
NOR2_X1 _20046_ ( .A1(_10033_ ), .A2(_03075_ ), .ZN(_05263_ ) );
NOR2_X1 _20047_ ( .A1(_05263_ ), .A2(\u_lsu.pmem[1127] ), .ZN(_05264_ ) );
AOI211_X1 _20048_ ( .A(fanout_net_68 ), .B(_05264_ ), .C1(_04216_ ), .C2(_05263_ ), .ZN(_01981_ ) );
NAND4_X1 _20049_ ( .A1(_05199_ ), .A2(_09925_ ), .A3(_05238_ ), .A4(_10930_ ), .ZN(_05265_ ) );
OAI21_X1 _20050_ ( .A(\u_lsu.pmem[1126] ), .B1(_05131_ ), .B2(_03076_ ), .ZN(_05266_ ) );
AOI21_X1 _20051_ ( .A(fanout_net_68 ), .B1(_05265_ ), .B2(_05266_ ), .ZN(_01982_ ) );
NAND4_X1 _20052_ ( .A1(_05199_ ), .A2(_09928_ ), .A3(_05238_ ), .A4(_10930_ ), .ZN(_05267_ ) );
OAI21_X1 _20053_ ( .A(\u_lsu.pmem[1125] ), .B1(_05131_ ), .B2(_03076_ ), .ZN(_05268_ ) );
AOI21_X1 _20054_ ( .A(fanout_net_68 ), .B1(_05267_ ), .B2(_05268_ ), .ZN(_01983_ ) );
NAND4_X1 _20055_ ( .A1(_05199_ ), .A2(_09931_ ), .A3(_05238_ ), .A4(_10930_ ), .ZN(_05269_ ) );
OAI21_X1 _20056_ ( .A(\u_lsu.pmem[1124] ), .B1(_05131_ ), .B2(_03075_ ), .ZN(_05270_ ) );
AOI21_X1 _20057_ ( .A(fanout_net_68 ), .B1(_05269_ ), .B2(_05270_ ), .ZN(_01984_ ) );
NAND4_X1 _20058_ ( .A1(_05199_ ), .A2(_03091_ ), .A3(_05238_ ), .A4(_10930_ ), .ZN(_05271_ ) );
OAI21_X1 _20059_ ( .A(\u_lsu.pmem[1123] ), .B1(_05131_ ), .B2(_03075_ ), .ZN(_05272_ ) );
AOI21_X1 _20060_ ( .A(fanout_net_68 ), .B1(_05271_ ), .B2(_05272_ ), .ZN(_01985_ ) );
NAND4_X1 _20061_ ( .A1(_05199_ ), .A2(_09938_ ), .A3(_05238_ ), .A4(_10930_ ), .ZN(_05273_ ) );
OAI21_X1 _20062_ ( .A(\u_lsu.pmem[1122] ), .B1(_05131_ ), .B2(_03075_ ), .ZN(_05274_ ) );
AOI21_X1 _20063_ ( .A(fanout_net_68 ), .B1(_05273_ ), .B2(_05274_ ), .ZN(_01986_ ) );
NAND4_X1 _20064_ ( .A1(_05199_ ), .A2(_03143_ ), .A3(_05238_ ), .A4(_10930_ ), .ZN(_05275_ ) );
OAI21_X1 _20065_ ( .A(\u_lsu.pmem[1121] ), .B1(_05131_ ), .B2(_03075_ ), .ZN(_05276_ ) );
AOI21_X1 _20066_ ( .A(fanout_net_68 ), .B1(_05275_ ), .B2(_05276_ ), .ZN(_01987_ ) );
BUF_X4 _20067_ ( .A(_10063_ ), .Z(_05277_ ) );
NAND4_X1 _20068_ ( .A1(_10088_ ), .A2(_05277_ ), .A3(_04658_ ), .A4(_05223_ ), .ZN(_05278_ ) );
OAI21_X1 _20069_ ( .A(\u_lsu.pmem[4066] ), .B1(_10068_ ), .B2(_04671_ ), .ZN(_05279_ ) );
AOI21_X1 _20070_ ( .A(fanout_net_68 ), .B1(_05278_ ), .B2(_05279_ ), .ZN(_01988_ ) );
NAND4_X1 _20071_ ( .A1(_05199_ ), .A2(_09944_ ), .A3(_05238_ ), .A4(_10930_ ), .ZN(_05280_ ) );
OAI21_X1 _20072_ ( .A(\u_lsu.pmem[1120] ), .B1(_05131_ ), .B2(_03075_ ), .ZN(_05281_ ) );
AOI21_X1 _20073_ ( .A(fanout_net_68 ), .B1(_05280_ ), .B2(_05281_ ), .ZN(_01989_ ) );
NOR2_X1 _20074_ ( .A1(_10033_ ), .A2(_03100_ ), .ZN(_05282_ ) );
NOR2_X1 _20075_ ( .A1(_05282_ ), .A2(\u_lsu.pmem[1095] ), .ZN(_05283_ ) );
AOI211_X1 _20076_ ( .A(fanout_net_68 ), .B(_05283_ ), .C1(_09567_ ), .C2(_05282_ ), .ZN(_01990_ ) );
NAND4_X1 _20077_ ( .A1(_05199_ ), .A2(_09957_ ), .A3(_09876_ ), .A4(_05011_ ), .ZN(_05284_ ) );
BUF_X4 _20078_ ( .A(_09472_ ), .Z(_05285_ ) );
OAI21_X1 _20079_ ( .A(\u_lsu.pmem[1094] ), .B1(_05285_ ), .B2(_03101_ ), .ZN(_05286_ ) );
AOI21_X1 _20080_ ( .A(fanout_net_68 ), .B1(_05284_ ), .B2(_05286_ ), .ZN(_01991_ ) );
NAND4_X1 _20081_ ( .A1(_05199_ ), .A2(_09961_ ), .A3(_09876_ ), .A4(_05011_ ), .ZN(_05287_ ) );
OAI21_X1 _20082_ ( .A(\u_lsu.pmem[1093] ), .B1(_05285_ ), .B2(_03101_ ), .ZN(_05288_ ) );
AOI21_X1 _20083_ ( .A(fanout_net_68 ), .B1(_05287_ ), .B2(_05288_ ), .ZN(_01992_ ) );
BUF_X4 _20084_ ( .A(_10036_ ), .Z(_05289_ ) );
NAND4_X1 _20085_ ( .A1(_05289_ ), .A2(_09966_ ), .A3(_09876_ ), .A4(_05011_ ), .ZN(_05290_ ) );
OAI21_X1 _20086_ ( .A(\u_lsu.pmem[1092] ), .B1(_05285_ ), .B2(_03100_ ), .ZN(_05291_ ) );
AOI21_X1 _20087_ ( .A(fanout_net_68 ), .B1(_05290_ ), .B2(_05291_ ), .ZN(_01993_ ) );
NAND4_X1 _20088_ ( .A1(_05289_ ), .A2(_09970_ ), .A3(_09876_ ), .A4(_05011_ ), .ZN(_05292_ ) );
OAI21_X1 _20089_ ( .A(\u_lsu.pmem[1091] ), .B1(_05285_ ), .B2(_03100_ ), .ZN(_05293_ ) );
AOI21_X1 _20090_ ( .A(fanout_net_68 ), .B1(_05292_ ), .B2(_05293_ ), .ZN(_01994_ ) );
NAND4_X1 _20091_ ( .A1(_05289_ ), .A2(_09974_ ), .A3(_09876_ ), .A4(_05011_ ), .ZN(_05294_ ) );
OAI21_X1 _20092_ ( .A(\u_lsu.pmem[1090] ), .B1(_05285_ ), .B2(_03100_ ), .ZN(_05295_ ) );
AOI21_X1 _20093_ ( .A(fanout_net_68 ), .B1(_05294_ ), .B2(_05295_ ), .ZN(_01995_ ) );
NAND4_X1 _20094_ ( .A1(_05289_ ), .A2(_09978_ ), .A3(_09876_ ), .A4(_05011_ ), .ZN(_05296_ ) );
OAI21_X1 _20095_ ( .A(\u_lsu.pmem[1089] ), .B1(_05285_ ), .B2(_03100_ ), .ZN(_05297_ ) );
AOI21_X1 _20096_ ( .A(fanout_net_68 ), .B1(_05296_ ), .B2(_05297_ ), .ZN(_01996_ ) );
NAND4_X1 _20097_ ( .A1(_05289_ ), .A2(_09982_ ), .A3(_09876_ ), .A4(_05011_ ), .ZN(_05298_ ) );
OAI21_X1 _20098_ ( .A(\u_lsu.pmem[1088] ), .B1(_05285_ ), .B2(_03100_ ), .ZN(_05299_ ) );
AOI21_X1 _20099_ ( .A(fanout_net_68 ), .B1(_05298_ ), .B2(_05299_ ), .ZN(_01997_ ) );
BUF_X4 _20100_ ( .A(_05166_ ), .Z(_05300_ ) );
NAND4_X1 _20101_ ( .A1(_09987_ ), .A2(_05277_ ), .A3(_05238_ ), .A4(_05300_ ), .ZN(_05301_ ) );
OAI21_X1 _20102_ ( .A(\u_lsu.pmem[1063] ), .B1(_05285_ ), .B2(_03127_ ), .ZN(_05302_ ) );
AOI21_X1 _20103_ ( .A(fanout_net_68 ), .B1(_05301_ ), .B2(_05302_ ), .ZN(_01998_ ) );
NAND4_X1 _20104_ ( .A1(_10094_ ), .A2(_05277_ ), .A3(_04658_ ), .A4(_05300_ ), .ZN(_05303_ ) );
OAI21_X1 _20105_ ( .A(\u_lsu.pmem[4065] ), .B1(_10068_ ), .B2(_04671_ ), .ZN(_05304_ ) );
AOI21_X1 _20106_ ( .A(fanout_net_68 ), .B1(_05303_ ), .B2(_05304_ ), .ZN(_01999_ ) );
BUF_X4 _20107_ ( .A(_05181_ ), .Z(_05305_ ) );
NAND4_X1 _20108_ ( .A1(_09994_ ), .A2(_05277_ ), .A3(_05305_ ), .A4(_05300_ ), .ZN(_05306_ ) );
OAI21_X1 _20109_ ( .A(\u_lsu.pmem[1062] ), .B1(_05285_ ), .B2(_03127_ ), .ZN(_05307_ ) );
AOI21_X1 _20110_ ( .A(fanout_net_68 ), .B1(_05306_ ), .B2(_05307_ ), .ZN(_02000_ ) );
NAND4_X1 _20111_ ( .A1(_09997_ ), .A2(_05277_ ), .A3(_05305_ ), .A4(_05300_ ), .ZN(_05308_ ) );
OAI21_X1 _20112_ ( .A(\u_lsu.pmem[1061] ), .B1(_05285_ ), .B2(_03126_ ), .ZN(_05309_ ) );
AOI21_X1 _20113_ ( .A(fanout_net_68 ), .B1(_05308_ ), .B2(_05309_ ), .ZN(_02001_ ) );
NAND4_X1 _20114_ ( .A1(_05289_ ), .A2(_09931_ ), .A3(_05305_ ), .A4(_10988_ ), .ZN(_05310_ ) );
OAI21_X1 _20115_ ( .A(\u_lsu.pmem[1060] ), .B1(_10785_ ), .B2(_03126_ ), .ZN(_05311_ ) );
AOI21_X1 _20116_ ( .A(fanout_net_69 ), .B1(_05310_ ), .B2(_05311_ ), .ZN(_02002_ ) );
NAND4_X1 _20117_ ( .A1(_05289_ ), .A2(_09934_ ), .A3(_05305_ ), .A4(_10988_ ), .ZN(_05312_ ) );
OAI21_X1 _20118_ ( .A(\u_lsu.pmem[1059] ), .B1(_10785_ ), .B2(_03126_ ), .ZN(_05313_ ) );
AOI21_X1 _20119_ ( .A(fanout_net_69 ), .B1(_05312_ ), .B2(_05313_ ), .ZN(_02003_ ) );
NAND4_X1 _20120_ ( .A1(_05289_ ), .A2(_09938_ ), .A3(_05305_ ), .A4(_10988_ ), .ZN(_05314_ ) );
OAI21_X1 _20121_ ( .A(\u_lsu.pmem[1058] ), .B1(_10785_ ), .B2(_03126_ ), .ZN(_05315_ ) );
AOI21_X1 _20122_ ( .A(fanout_net_69 ), .B1(_05314_ ), .B2(_05315_ ), .ZN(_02004_ ) );
NAND4_X1 _20123_ ( .A1(_05289_ ), .A2(_09941_ ), .A3(_05305_ ), .A4(_10988_ ), .ZN(_05316_ ) );
OAI21_X1 _20124_ ( .A(\u_lsu.pmem[1057] ), .B1(_10785_ ), .B2(_03126_ ), .ZN(_05317_ ) );
AOI21_X1 _20125_ ( .A(fanout_net_69 ), .B1(_05316_ ), .B2(_05317_ ), .ZN(_02005_ ) );
NAND4_X1 _20126_ ( .A1(_10021_ ), .A2(_05277_ ), .A3(_05305_ ), .A4(_05300_ ), .ZN(_05318_ ) );
OAI21_X1 _20127_ ( .A(\u_lsu.pmem[1056] ), .B1(_10785_ ), .B2(_03126_ ), .ZN(_05319_ ) );
AOI21_X1 _20128_ ( .A(fanout_net_69 ), .B1(_05318_ ), .B2(_05319_ ), .ZN(_02006_ ) );
NAND4_X1 _20129_ ( .A1(_09700_ ), .A2(_09603_ ), .A3(_10071_ ), .A4(_03151_ ), .ZN(_05320_ ) );
BUF_X4 _20130_ ( .A(_10041_ ), .Z(_05321_ ) );
OAI21_X1 _20131_ ( .A(\u_lsu.pmem[1031] ), .B1(_03155_ ), .B2(_05321_ ), .ZN(_05322_ ) );
AOI21_X1 _20132_ ( .A(fanout_net_69 ), .B1(_05320_ ), .B2(_05322_ ), .ZN(_02007_ ) );
NAND3_X1 _20133_ ( .A1(_05008_ ), .A2(_11145_ ), .A3(_03151_ ), .ZN(_05323_ ) );
OAI21_X1 _20134_ ( .A(\u_lsu.pmem[1030] ), .B1(_03155_ ), .B2(_05321_ ), .ZN(_05324_ ) );
AOI21_X1 _20135_ ( .A(fanout_net_69 ), .B1(_05323_ ), .B2(_05324_ ), .ZN(_02008_ ) );
NAND3_X1 _20136_ ( .A1(_05008_ ), .A2(_11148_ ), .A3(_03151_ ), .ZN(_05325_ ) );
OAI21_X1 _20137_ ( .A(\u_lsu.pmem[1029] ), .B1(_03155_ ), .B2(_05321_ ), .ZN(_05326_ ) );
AOI21_X1 _20138_ ( .A(fanout_net_69 ), .B1(_05325_ ), .B2(_05326_ ), .ZN(_02009_ ) );
NAND4_X1 _20139_ ( .A1(_10098_ ), .A2(_05277_ ), .A3(_04658_ ), .A4(_05300_ ), .ZN(_05327_ ) );
OAI21_X1 _20140_ ( .A(\u_lsu.pmem[4064] ), .B1(_10068_ ), .B2(_05321_ ), .ZN(_05328_ ) );
AOI21_X1 _20141_ ( .A(fanout_net_69 ), .B1(_05327_ ), .B2(_05328_ ), .ZN(_02010_ ) );
NAND3_X1 _20142_ ( .A1(_05008_ ), .A2(_03084_ ), .A3(_03151_ ), .ZN(_05329_ ) );
OAI21_X1 _20143_ ( .A(\u_lsu.pmem[1028] ), .B1(_03155_ ), .B2(_05321_ ), .ZN(_05330_ ) );
AOI21_X1 _20144_ ( .A(fanout_net_69 ), .B1(_05329_ ), .B2(_05330_ ), .ZN(_02011_ ) );
NAND3_X1 _20145_ ( .A1(_05008_ ), .A2(_11155_ ), .A3(_03151_ ), .ZN(_05331_ ) );
OAI21_X1 _20146_ ( .A(\u_lsu.pmem[1027] ), .B1(_03155_ ), .B2(_05321_ ), .ZN(_05332_ ) );
AOI21_X1 _20147_ ( .A(fanout_net_69 ), .B1(_05331_ ), .B2(_05332_ ), .ZN(_02012_ ) );
NAND4_X1 _20148_ ( .A1(_11021_ ), .A2(_04914_ ), .A3(_05305_ ), .A4(_05300_ ), .ZN(_05333_ ) );
OAI21_X1 _20149_ ( .A(\u_lsu.pmem[1026] ), .B1(_03155_ ), .B2(_05321_ ), .ZN(_05334_ ) );
AOI21_X1 _20150_ ( .A(fanout_net_69 ), .B1(_05333_ ), .B2(_05334_ ), .ZN(_02013_ ) );
NAND3_X1 _20151_ ( .A1(_05008_ ), .A2(_11163_ ), .A3(_03151_ ), .ZN(_05335_ ) );
OAI21_X1 _20152_ ( .A(\u_lsu.pmem[1025] ), .B1(_03155_ ), .B2(_05321_ ), .ZN(_05336_ ) );
AOI21_X1 _20153_ ( .A(fanout_net_69 ), .B1(_05335_ ), .B2(_05336_ ), .ZN(_02014_ ) );
NAND3_X1 _20154_ ( .A1(_05008_ ), .A2(_03203_ ), .A3(_03151_ ), .ZN(_05337_ ) );
OAI21_X1 _20155_ ( .A(\u_lsu.pmem[1024] ), .B1(_03155_ ), .B2(_05321_ ), .ZN(_05338_ ) );
AOI21_X1 _20156_ ( .A(fanout_net_69 ), .B1(_05337_ ), .B2(_05338_ ), .ZN(_02015_ ) );
NAND4_X1 _20157_ ( .A1(_05289_ ), .A2(_09674_ ), .A3(_04928_ ), .A4(_11030_ ), .ZN(_05339_ ) );
OAI21_X1 _20158_ ( .A(\u_lsu.pmem[999] ), .B1(_03171_ ), .B2(_05221_ ), .ZN(_05340_ ) );
AOI21_X1 _20159_ ( .A(fanout_net_69 ), .B1(_05339_ ), .B2(_05340_ ), .ZN(_02016_ ) );
NAND4_X1 _20160_ ( .A1(_10062_ ), .A2(_04914_ ), .A3(_05305_ ), .A4(_05300_ ), .ZN(_05341_ ) );
OAI21_X1 _20161_ ( .A(\u_lsu.pmem[998] ), .B1(_03171_ ), .B2(_05221_ ), .ZN(_05342_ ) );
AOI21_X1 _20162_ ( .A(fanout_net_69 ), .B1(_05341_ ), .B2(_05342_ ), .ZN(_02017_ ) );
NAND4_X1 _20163_ ( .A1(_10075_ ), .A2(_04914_ ), .A3(_05305_ ), .A4(_05300_ ), .ZN(_05343_ ) );
BUF_X4 _20164_ ( .A(_05046_ ), .Z(_05344_ ) );
OAI21_X1 _20165_ ( .A(\u_lsu.pmem[997] ), .B1(_03171_ ), .B2(_05344_ ), .ZN(_05345_ ) );
AOI21_X1 _20166_ ( .A(fanout_net_69 ), .B1(_05343_ ), .B2(_05345_ ), .ZN(_02018_ ) );
BUF_X4 _20167_ ( .A(_05181_ ), .Z(_05346_ ) );
NAND4_X1 _20168_ ( .A1(_10079_ ), .A2(_04914_ ), .A3(_05346_ ), .A4(_05300_ ), .ZN(_05347_ ) );
OAI21_X1 _20169_ ( .A(\u_lsu.pmem[996] ), .B1(_03171_ ), .B2(_05344_ ), .ZN(_05348_ ) );
AOI21_X1 _20170_ ( .A(fanout_net_69 ), .B1(_05347_ ), .B2(_05348_ ), .ZN(_02019_ ) );
BUF_X4 _20171_ ( .A(_05166_ ), .Z(_05349_ ) );
NAND4_X1 _20172_ ( .A1(_10084_ ), .A2(_04914_ ), .A3(_05346_ ), .A4(_05349_ ), .ZN(_05350_ ) );
OAI21_X1 _20173_ ( .A(\u_lsu.pmem[995] ), .B1(_03171_ ), .B2(_05344_ ), .ZN(_05351_ ) );
AOI21_X1 _20174_ ( .A(fanout_net_69 ), .B1(_05350_ ), .B2(_05351_ ), .ZN(_02020_ ) );
AND2_X1 _20175_ ( .A1(_10105_ ), .A2(_11011_ ), .ZN(_05352_ ) );
OAI21_X1 _20176_ ( .A(_09109_ ), .B1(_05352_ ), .B2(\u_lsu.pmem[4039] ), .ZN(_05353_ ) );
AOI21_X1 _20177_ ( .A(_05353_ ), .B1(_09568_ ), .B2(_05352_ ), .ZN(_02021_ ) );
NAND4_X1 _20178_ ( .A1(_10088_ ), .A2(_04914_ ), .A3(_05346_ ), .A4(_05349_ ), .ZN(_05354_ ) );
OAI21_X1 _20179_ ( .A(\u_lsu.pmem[994] ), .B1(_03171_ ), .B2(_05344_ ), .ZN(_05355_ ) );
AOI21_X1 _20180_ ( .A(fanout_net_69 ), .B1(_05354_ ), .B2(_05355_ ), .ZN(_02022_ ) );
NAND4_X1 _20181_ ( .A1(_10094_ ), .A2(_04914_ ), .A3(_05346_ ), .A4(_05349_ ), .ZN(_05356_ ) );
OAI21_X1 _20182_ ( .A(\u_lsu.pmem[993] ), .B1(_03171_ ), .B2(_05344_ ), .ZN(_05357_ ) );
AOI21_X1 _20183_ ( .A(fanout_net_69 ), .B1(_05356_ ), .B2(_05357_ ), .ZN(_02023_ ) );
BUF_X4 _20184_ ( .A(_04210_ ), .Z(_05358_ ) );
NAND4_X1 _20185_ ( .A1(_10098_ ), .A2(_05358_ ), .A3(_05346_ ), .A4(_05349_ ), .ZN(_05359_ ) );
OAI21_X1 _20186_ ( .A(\u_lsu.pmem[992] ), .B1(_03171_ ), .B2(_05344_ ), .ZN(_05360_ ) );
AOI21_X1 _20187_ ( .A(fanout_net_69 ), .B1(_05359_ ), .B2(_05360_ ), .ZN(_02024_ ) );
NAND4_X1 _20188_ ( .A1(_10037_ ), .A2(_09674_ ), .A3(_04928_ ), .A4(_11057_ ), .ZN(_05361_ ) );
OAI21_X1 _20189_ ( .A(\u_lsu.pmem[967] ), .B1(_03196_ ), .B2(_05344_ ), .ZN(_05362_ ) );
AOI21_X1 _20190_ ( .A(fanout_net_69 ), .B1(_05361_ ), .B2(_05362_ ), .ZN(_02025_ ) );
NAND4_X1 _20191_ ( .A1(_10117_ ), .A2(_05358_ ), .A3(_05346_ ), .A4(_05349_ ), .ZN(_05363_ ) );
OAI21_X1 _20192_ ( .A(\u_lsu.pmem[966] ), .B1(_03196_ ), .B2(_05344_ ), .ZN(_05364_ ) );
AOI21_X1 _20193_ ( .A(fanout_net_69 ), .B1(_05363_ ), .B2(_05364_ ), .ZN(_02026_ ) );
NAND4_X1 _20194_ ( .A1(_10121_ ), .A2(_05358_ ), .A3(_05346_ ), .A4(_05349_ ), .ZN(_05365_ ) );
OAI21_X1 _20195_ ( .A(\u_lsu.pmem[965] ), .B1(_03196_ ), .B2(_05344_ ), .ZN(_05366_ ) );
AOI21_X1 _20196_ ( .A(fanout_net_69 ), .B1(_05365_ ), .B2(_05366_ ), .ZN(_02027_ ) );
NAND4_X1 _20197_ ( .A1(_10125_ ), .A2(_05358_ ), .A3(_05346_ ), .A4(_05349_ ), .ZN(_05367_ ) );
OAI21_X1 _20198_ ( .A(\u_lsu.pmem[964] ), .B1(_03196_ ), .B2(_05344_ ), .ZN(_05368_ ) );
AOI21_X1 _20199_ ( .A(fanout_net_69 ), .B1(_05367_ ), .B2(_05368_ ), .ZN(_02028_ ) );
NAND4_X1 _20200_ ( .A1(_10131_ ), .A2(_05358_ ), .A3(_05346_ ), .A4(_05349_ ), .ZN(_05369_ ) );
BUF_X4 _20201_ ( .A(_05046_ ), .Z(_05370_ ) );
OAI21_X1 _20202_ ( .A(\u_lsu.pmem[963] ), .B1(_03196_ ), .B2(_05370_ ), .ZN(_05371_ ) );
AOI21_X1 _20203_ ( .A(fanout_net_69 ), .B1(_05369_ ), .B2(_05371_ ), .ZN(_02029_ ) );
NAND4_X1 _20204_ ( .A1(_10135_ ), .A2(_05358_ ), .A3(_05346_ ), .A4(_05349_ ), .ZN(_05372_ ) );
OAI21_X1 _20205_ ( .A(\u_lsu.pmem[962] ), .B1(_03196_ ), .B2(_05370_ ), .ZN(_05373_ ) );
AOI21_X1 _20206_ ( .A(fanout_net_69 ), .B1(_05372_ ), .B2(_05373_ ), .ZN(_02030_ ) );
BUF_X4 _20207_ ( .A(_05181_ ), .Z(_05374_ ) );
NAND4_X1 _20208_ ( .A1(_10138_ ), .A2(_05358_ ), .A3(_05374_ ), .A4(_05349_ ), .ZN(_05375_ ) );
OAI21_X1 _20209_ ( .A(\u_lsu.pmem[961] ), .B1(_03196_ ), .B2(_05370_ ), .ZN(_05376_ ) );
AOI21_X1 _20210_ ( .A(fanout_net_69 ), .B1(_05375_ ), .B2(_05376_ ), .ZN(_02031_ ) );
BUF_X4 _20211_ ( .A(_05166_ ), .Z(_05377_ ) );
NAND4_X1 _20212_ ( .A1(_10117_ ), .A2(_05277_ ), .A3(_04658_ ), .A4(_05377_ ), .ZN(_05378_ ) );
OAI21_X1 _20213_ ( .A(\u_lsu.pmem[4038] ), .B1(_10107_ ), .B2(_05321_ ), .ZN(_05379_ ) );
AOI21_X1 _20214_ ( .A(fanout_net_69 ), .B1(_05378_ ), .B2(_05379_ ), .ZN(_02032_ ) );
NAND4_X1 _20215_ ( .A1(_10144_ ), .A2(_05358_ ), .A3(_05374_ ), .A4(_05377_ ), .ZN(_05380_ ) );
OAI21_X1 _20216_ ( .A(\u_lsu.pmem[960] ), .B1(_03196_ ), .B2(_05370_ ), .ZN(_05381_ ) );
AOI21_X1 _20217_ ( .A(fanout_net_70 ), .B1(_05380_ ), .B2(_05381_ ), .ZN(_02033_ ) );
NAND4_X1 _20218_ ( .A1(_10148_ ), .A2(_05358_ ), .A3(_05374_ ), .A4(_05377_ ), .ZN(_05382_ ) );
OAI21_X1 _20219_ ( .A(\u_lsu.pmem[935] ), .B1(_03222_ ), .B2(_05370_ ), .ZN(_05383_ ) );
AOI21_X1 _20220_ ( .A(fanout_net_70 ), .B1(_05382_ ), .B2(_05383_ ), .ZN(_02034_ ) );
NAND4_X1 _20221_ ( .A1(_10156_ ), .A2(_05358_ ), .A3(_05374_ ), .A4(_05377_ ), .ZN(_05384_ ) );
OAI21_X1 _20222_ ( .A(\u_lsu.pmem[934] ), .B1(_03222_ ), .B2(_05370_ ), .ZN(_05385_ ) );
AOI21_X1 _20223_ ( .A(fanout_net_70 ), .B1(_05384_ ), .B2(_05385_ ), .ZN(_02035_ ) );
BUF_X4 _20224_ ( .A(_09883_ ), .Z(_05386_ ) );
NAND4_X1 _20225_ ( .A1(_10160_ ), .A2(_05386_ ), .A3(_05374_ ), .A4(_05377_ ), .ZN(_05387_ ) );
OAI21_X1 _20226_ ( .A(\u_lsu.pmem[933] ), .B1(_03222_ ), .B2(_05370_ ), .ZN(_05388_ ) );
AOI21_X1 _20227_ ( .A(fanout_net_70 ), .B1(_05387_ ), .B2(_05388_ ), .ZN(_02036_ ) );
NAND4_X1 _20228_ ( .A1(_10166_ ), .A2(_05386_ ), .A3(_05374_ ), .A4(_05377_ ), .ZN(_05389_ ) );
OAI21_X1 _20229_ ( .A(\u_lsu.pmem[932] ), .B1(_03222_ ), .B2(_05370_ ), .ZN(_05390_ ) );
AOI21_X1 _20230_ ( .A(fanout_net_70 ), .B1(_05389_ ), .B2(_05390_ ), .ZN(_02037_ ) );
NAND4_X1 _20231_ ( .A1(_10169_ ), .A2(_05386_ ), .A3(_05374_ ), .A4(_05377_ ), .ZN(_05391_ ) );
OAI21_X1 _20232_ ( .A(\u_lsu.pmem[931] ), .B1(_03222_ ), .B2(_05370_ ), .ZN(_05392_ ) );
AOI21_X1 _20233_ ( .A(fanout_net_70 ), .B1(_05391_ ), .B2(_05392_ ), .ZN(_02038_ ) );
NAND4_X1 _20234_ ( .A1(_10172_ ), .A2(_05386_ ), .A3(_05374_ ), .A4(_05377_ ), .ZN(_05393_ ) );
OAI21_X1 _20235_ ( .A(\u_lsu.pmem[930] ), .B1(_03222_ ), .B2(_05370_ ), .ZN(_05394_ ) );
AOI21_X1 _20236_ ( .A(fanout_net_70 ), .B1(_05393_ ), .B2(_05394_ ), .ZN(_02039_ ) );
NAND4_X1 _20237_ ( .A1(_10176_ ), .A2(_05386_ ), .A3(_05374_ ), .A4(_05377_ ), .ZN(_05395_ ) );
BUF_X4 _20238_ ( .A(_05046_ ), .Z(_05396_ ) );
OAI21_X1 _20239_ ( .A(\u_lsu.pmem[929] ), .B1(_03222_ ), .B2(_05396_ ), .ZN(_05397_ ) );
AOI21_X1 _20240_ ( .A(fanout_net_70 ), .B1(_05395_ ), .B2(_05397_ ), .ZN(_02040_ ) );
NAND4_X1 _20241_ ( .A1(_10037_ ), .A2(_09944_ ), .A3(_05374_ ), .A4(_11086_ ), .ZN(_05398_ ) );
OAI21_X1 _20242_ ( .A(\u_lsu.pmem[928] ), .B1(_03222_ ), .B2(_05396_ ), .ZN(_05399_ ) );
AOI21_X1 _20243_ ( .A(fanout_net_70 ), .B1(_05398_ ), .B2(_05399_ ), .ZN(_02041_ ) );
OAI21_X1 _20244_ ( .A(\u_lsu.pmem[903] ), .B1(_03246_ ), .B2(_05247_ ), .ZN(_05400_ ) );
BUF_X4 _20245_ ( .A(_09455_ ), .Z(_05401_ ) );
NAND4_X1 _20246_ ( .A1(_11112_ ), .A2(_08582_ ), .A3(_05401_ ), .A4(_05257_ ), .ZN(_05402_ ) );
AOI21_X1 _20247_ ( .A(fanout_net_70 ), .B1(_05400_ ), .B2(_05402_ ), .ZN(_02042_ ) );
NAND4_X1 _20248_ ( .A1(_10121_ ), .A2(_05277_ ), .A3(_04658_ ), .A4(_05377_ ), .ZN(_05403_ ) );
OAI21_X1 _20249_ ( .A(\u_lsu.pmem[4037] ), .B1(_10107_ ), .B2(_10110_ ), .ZN(_05404_ ) );
AOI21_X1 _20250_ ( .A(fanout_net_70 ), .B1(_05403_ ), .B2(_05404_ ), .ZN(_02043_ ) );
OAI21_X1 _20251_ ( .A(\u_lsu.pmem[902] ), .B1(_03246_ ), .B2(_05247_ ), .ZN(_05405_ ) );
NAND4_X1 _20252_ ( .A1(_11112_ ), .A2(_09575_ ), .A3(_05401_ ), .A4(_05257_ ), .ZN(_05406_ ) );
AOI21_X1 _20253_ ( .A(fanout_net_70 ), .B1(_05405_ ), .B2(_05406_ ), .ZN(_02044_ ) );
OAI21_X1 _20254_ ( .A(\u_lsu.pmem[901] ), .B1(_03245_ ), .B2(_05247_ ), .ZN(_05407_ ) );
NAND4_X1 _20255_ ( .A1(_11112_ ), .A2(_09582_ ), .A3(_05401_ ), .A4(_05257_ ), .ZN(_05408_ ) );
AOI21_X1 _20256_ ( .A(fanout_net_70 ), .B1(_05407_ ), .B2(_05408_ ), .ZN(_02045_ ) );
OAI21_X1 _20257_ ( .A(\u_lsu.pmem[900] ), .B1(_03245_ ), .B2(_05247_ ), .ZN(_05409_ ) );
NAND4_X1 _20258_ ( .A1(_11112_ ), .A2(_08605_ ), .A3(_05401_ ), .A4(_05257_ ), .ZN(_05410_ ) );
AOI21_X1 _20259_ ( .A(fanout_net_70 ), .B1(_05409_ ), .B2(_05410_ ), .ZN(_02046_ ) );
BUF_X4 _20260_ ( .A(_10720_ ), .Z(_05411_ ) );
OAI21_X1 _20261_ ( .A(\u_lsu.pmem[899] ), .B1(_03245_ ), .B2(_05411_ ), .ZN(_05412_ ) );
NAND4_X1 _20262_ ( .A1(_11112_ ), .A2(_09519_ ), .A3(_05401_ ), .A4(_05257_ ), .ZN(_05413_ ) );
AOI21_X1 _20263_ ( .A(fanout_net_70 ), .B1(_05412_ ), .B2(_05413_ ), .ZN(_02047_ ) );
OAI21_X1 _20264_ ( .A(\u_lsu.pmem[898] ), .B1(_03245_ ), .B2(_05411_ ), .ZN(_05414_ ) );
NAND4_X1 _20265_ ( .A1(_09874_ ), .A2(_04585_ ), .A3(_05401_ ), .A4(_05257_ ), .ZN(_05415_ ) );
AOI21_X1 _20266_ ( .A(fanout_net_70 ), .B1(_05414_ ), .B2(_05415_ ), .ZN(_02048_ ) );
OAI21_X1 _20267_ ( .A(\u_lsu.pmem[897] ), .B1(_03245_ ), .B2(_05411_ ), .ZN(_05416_ ) );
NAND4_X1 _20268_ ( .A1(_11112_ ), .A2(_09543_ ), .A3(_05401_ ), .A4(_05257_ ), .ZN(_05417_ ) );
AOI21_X1 _20269_ ( .A(fanout_net_70 ), .B1(_05416_ ), .B2(_05417_ ), .ZN(_02049_ ) );
OAI21_X1 _20270_ ( .A(\u_lsu.pmem[896] ), .B1(_03245_ ), .B2(_05411_ ), .ZN(_05418_ ) );
NAND4_X1 _20271_ ( .A1(_11112_ ), .A2(_09547_ ), .A3(_05401_ ), .A4(_04008_ ), .ZN(_05419_ ) );
AOI21_X1 _20272_ ( .A(fanout_net_70 ), .B1(_05418_ ), .B2(_05419_ ), .ZN(_02050_ ) );
NAND3_X1 _20273_ ( .A1(_05008_ ), .A2(_11138_ ), .A3(_03276_ ), .ZN(_05420_ ) );
OAI21_X1 _20274_ ( .A(\u_lsu.pmem[871] ), .B1(_03273_ ), .B2(_05396_ ), .ZN(_05421_ ) );
AOI21_X1 _20275_ ( .A(fanout_net_70 ), .B1(_05420_ ), .B2(_05421_ ), .ZN(_02051_ ) );
BUF_X4 _20276_ ( .A(_09641_ ), .Z(_05422_ ) );
NAND3_X1 _20277_ ( .A1(_05422_ ), .A2(_11145_ ), .A3(_03276_ ), .ZN(_05423_ ) );
OAI21_X1 _20278_ ( .A(\u_lsu.pmem[870] ), .B1(_03273_ ), .B2(_05396_ ), .ZN(_05424_ ) );
AOI21_X1 _20279_ ( .A(fanout_net_70 ), .B1(_05423_ ), .B2(_05424_ ), .ZN(_02052_ ) );
NAND3_X1 _20280_ ( .A1(_05422_ ), .A2(_11148_ ), .A3(_03276_ ), .ZN(_05425_ ) );
OAI21_X1 _20281_ ( .A(\u_lsu.pmem[869] ), .B1(_03273_ ), .B2(_05396_ ), .ZN(_05426_ ) );
AOI21_X1 _20282_ ( .A(fanout_net_70 ), .B1(_05425_ ), .B2(_05426_ ), .ZN(_02053_ ) );
BUF_X4 _20283_ ( .A(_10578_ ), .Z(_05427_ ) );
BUF_X4 _20284_ ( .A(_05166_ ), .Z(_05428_ ) );
NAND4_X1 _20285_ ( .A1(_10125_ ), .A2(_05277_ ), .A3(_05427_ ), .A4(_05428_ ), .ZN(_05429_ ) );
OAI21_X1 _20286_ ( .A(\u_lsu.pmem[4036] ), .B1(_10106_ ), .B2(_10110_ ), .ZN(_05430_ ) );
AOI21_X1 _20287_ ( .A(fanout_net_70 ), .B1(_05429_ ), .B2(_05430_ ), .ZN(_02054_ ) );
NAND3_X1 _20288_ ( .A1(_05422_ ), .A2(_03084_ ), .A3(_03276_ ), .ZN(_05431_ ) );
OAI21_X1 _20289_ ( .A(\u_lsu.pmem[868] ), .B1(_03273_ ), .B2(_05396_ ), .ZN(_05432_ ) );
AOI21_X1 _20290_ ( .A(fanout_net_70 ), .B1(_05431_ ), .B2(_05432_ ), .ZN(_02055_ ) );
NAND3_X1 _20291_ ( .A1(_05422_ ), .A2(_11155_ ), .A3(_03276_ ), .ZN(_05433_ ) );
OAI21_X1 _20292_ ( .A(\u_lsu.pmem[867] ), .B1(_03273_ ), .B2(_05396_ ), .ZN(_05434_ ) );
AOI21_X1 _20293_ ( .A(fanout_net_70 ), .B1(_05433_ ), .B2(_05434_ ), .ZN(_02056_ ) );
NAND3_X1 _20294_ ( .A1(_05422_ ), .A2(_03145_ ), .A3(_03276_ ), .ZN(_05435_ ) );
OAI21_X1 _20295_ ( .A(\u_lsu.pmem[866] ), .B1(_03273_ ), .B2(_05396_ ), .ZN(_05436_ ) );
AOI21_X1 _20296_ ( .A(fanout_net_70 ), .B1(_05435_ ), .B2(_05436_ ), .ZN(_02057_ ) );
NAND3_X1 _20297_ ( .A1(_05422_ ), .A2(_11163_ ), .A3(_03276_ ), .ZN(_05437_ ) );
OAI21_X1 _20298_ ( .A(\u_lsu.pmem[865] ), .B1(_03273_ ), .B2(_05396_ ), .ZN(_05438_ ) );
AOI21_X1 _20299_ ( .A(fanout_net_70 ), .B1(_05437_ ), .B2(_05438_ ), .ZN(_02058_ ) );
NAND3_X1 _20300_ ( .A1(_05422_ ), .A2(_03203_ ), .A3(_03276_ ), .ZN(_05439_ ) );
OAI21_X1 _20301_ ( .A(\u_lsu.pmem[864] ), .B1(_03273_ ), .B2(_05396_ ), .ZN(_05440_ ) );
AOI21_X1 _20302_ ( .A(fanout_net_70 ), .B1(_05439_ ), .B2(_05440_ ), .ZN(_02059_ ) );
NAND3_X1 _20303_ ( .A1(_05422_ ), .A2(_11138_ ), .A3(_03297_ ), .ZN(_05441_ ) );
BUF_X4 _20304_ ( .A(_05046_ ), .Z(_05442_ ) );
OAI21_X1 _20305_ ( .A(\u_lsu.pmem[839] ), .B1(_03295_ ), .B2(_05442_ ), .ZN(_05443_ ) );
AOI21_X1 _20306_ ( .A(fanout_net_70 ), .B1(_05441_ ), .B2(_05443_ ), .ZN(_02060_ ) );
NAND3_X1 _20307_ ( .A1(_05422_ ), .A2(_11145_ ), .A3(_03297_ ), .ZN(_05444_ ) );
OAI21_X1 _20308_ ( .A(\u_lsu.pmem[838] ), .B1(_03295_ ), .B2(_05442_ ), .ZN(_05445_ ) );
AOI21_X1 _20309_ ( .A(fanout_net_70 ), .B1(_05444_ ), .B2(_05445_ ), .ZN(_02061_ ) );
NAND3_X1 _20310_ ( .A1(_05422_ ), .A2(_11148_ ), .A3(_03297_ ), .ZN(_05446_ ) );
OAI21_X1 _20311_ ( .A(\u_lsu.pmem[837] ), .B1(_03295_ ), .B2(_05442_ ), .ZN(_05447_ ) );
AOI21_X1 _20312_ ( .A(fanout_net_70 ), .B1(_05446_ ), .B2(_05447_ ), .ZN(_02062_ ) );
BUF_X4 _20313_ ( .A(_09641_ ), .Z(_05448_ ) );
NAND3_X1 _20314_ ( .A1(_05448_ ), .A2(_03084_ ), .A3(_03297_ ), .ZN(_05449_ ) );
OAI21_X1 _20315_ ( .A(\u_lsu.pmem[836] ), .B1(_03295_ ), .B2(_05442_ ), .ZN(_05450_ ) );
AOI21_X1 _20316_ ( .A(fanout_net_71 ), .B1(_05449_ ), .B2(_05450_ ), .ZN(_02063_ ) );
NAND3_X1 _20317_ ( .A1(_05448_ ), .A2(_11155_ ), .A3(_03297_ ), .ZN(_05451_ ) );
OAI21_X1 _20318_ ( .A(\u_lsu.pmem[835] ), .B1(_03295_ ), .B2(_05442_ ), .ZN(_05452_ ) );
AOI21_X1 _20319_ ( .A(fanout_net_71 ), .B1(_05451_ ), .B2(_05452_ ), .ZN(_02064_ ) );
BUF_X4 _20320_ ( .A(_10063_ ), .Z(_05453_ ) );
NAND4_X1 _20321_ ( .A1(_10131_ ), .A2(_05453_ ), .A3(_05427_ ), .A4(_05428_ ), .ZN(_05454_ ) );
OAI21_X1 _20322_ ( .A(\u_lsu.pmem[4035] ), .B1(_10106_ ), .B2(_10110_ ), .ZN(_05455_ ) );
AOI21_X1 _20323_ ( .A(fanout_net_71 ), .B1(_05454_ ), .B2(_05455_ ), .ZN(_02065_ ) );
NAND3_X1 _20324_ ( .A1(_05448_ ), .A2(_11158_ ), .A3(_03297_ ), .ZN(_05456_ ) );
OAI21_X1 _20325_ ( .A(\u_lsu.pmem[834] ), .B1(_03295_ ), .B2(_05442_ ), .ZN(_05457_ ) );
AOI21_X1 _20326_ ( .A(fanout_net_71 ), .B1(_05456_ ), .B2(_05457_ ), .ZN(_02066_ ) );
NAND3_X1 _20327_ ( .A1(_05448_ ), .A2(_11163_ ), .A3(_03297_ ), .ZN(_05458_ ) );
OAI21_X1 _20328_ ( .A(\u_lsu.pmem[833] ), .B1(_03295_ ), .B2(_05442_ ), .ZN(_05459_ ) );
AOI21_X1 _20329_ ( .A(fanout_net_71 ), .B1(_05458_ ), .B2(_05459_ ), .ZN(_02067_ ) );
NAND3_X1 _20330_ ( .A1(_05448_ ), .A2(_03203_ ), .A3(_03297_ ), .ZN(_05460_ ) );
OAI21_X1 _20331_ ( .A(\u_lsu.pmem[832] ), .B1(_03295_ ), .B2(_05442_ ), .ZN(_05461_ ) );
AOI21_X1 _20332_ ( .A(fanout_net_71 ), .B1(_05460_ ), .B2(_05461_ ), .ZN(_02068_ ) );
BUF_X4 _20333_ ( .A(_05181_ ), .Z(_05462_ ) );
NAND4_X1 _20334_ ( .A1(_10250_ ), .A2(_05386_ ), .A3(_05462_ ), .A4(_05428_ ), .ZN(_05463_ ) );
OAI21_X1 _20335_ ( .A(\u_lsu.pmem[807] ), .B1(_03335_ ), .B2(_05442_ ), .ZN(_05464_ ) );
AOI21_X1 _20336_ ( .A(fanout_net_71 ), .B1(_05463_ ), .B2(_05464_ ), .ZN(_02069_ ) );
NAND4_X1 _20337_ ( .A1(_10263_ ), .A2(_05386_ ), .A3(_05462_ ), .A4(_05428_ ), .ZN(_05465_ ) );
OAI21_X1 _20338_ ( .A(\u_lsu.pmem[806] ), .B1(_03335_ ), .B2(_05442_ ), .ZN(_05466_ ) );
AOI21_X1 _20339_ ( .A(fanout_net_71 ), .B1(_05465_ ), .B2(_05466_ ), .ZN(_02070_ ) );
NAND4_X1 _20340_ ( .A1(_10267_ ), .A2(_05386_ ), .A3(_05462_ ), .A4(_05428_ ), .ZN(_05467_ ) );
BUF_X4 _20341_ ( .A(_05046_ ), .Z(_05468_ ) );
OAI21_X1 _20342_ ( .A(\u_lsu.pmem[805] ), .B1(_03335_ ), .B2(_05468_ ), .ZN(_05469_ ) );
AOI21_X1 _20343_ ( .A(fanout_net_71 ), .B1(_05467_ ), .B2(_05469_ ), .ZN(_02071_ ) );
NOR2_X2 _20344_ ( .A1(_03321_ ), .A2(_09635_ ), .ZN(_05470_ ) );
OAI21_X1 _20345_ ( .A(_09109_ ), .B1(_05470_ ), .B2(\u_lsu.pmem[804] ), .ZN(_05471_ ) );
AOI21_X1 _20346_ ( .A(_05471_ ), .B1(_09149_ ), .B2(_05470_ ), .ZN(_02072_ ) );
NAND3_X1 _20347_ ( .A1(_05448_ ), .A2(_11155_ ), .A3(_03320_ ), .ZN(_05472_ ) );
OAI21_X1 _20348_ ( .A(\u_lsu.pmem[803] ), .B1(_03335_ ), .B2(_05468_ ), .ZN(_05473_ ) );
AOI21_X1 _20349_ ( .A(fanout_net_71 ), .B1(_05472_ ), .B2(_05473_ ), .ZN(_02073_ ) );
NAND3_X1 _20350_ ( .A1(_05448_ ), .A2(_11158_ ), .A3(_03320_ ), .ZN(_05474_ ) );
OAI21_X1 _20351_ ( .A(\u_lsu.pmem[802] ), .B1(_03335_ ), .B2(_05468_ ), .ZN(_05475_ ) );
AOI21_X1 _20352_ ( .A(fanout_net_71 ), .B1(_05474_ ), .B2(_05475_ ), .ZN(_02074_ ) );
NAND3_X1 _20353_ ( .A1(_05448_ ), .A2(_11163_ ), .A3(_03320_ ), .ZN(_05476_ ) );
OAI21_X1 _20354_ ( .A(\u_lsu.pmem[801] ), .B1(_03335_ ), .B2(_05468_ ), .ZN(_05477_ ) );
AOI21_X1 _20355_ ( .A(fanout_net_71 ), .B1(_05476_ ), .B2(_05477_ ), .ZN(_02075_ ) );
NAND4_X1 _20356_ ( .A1(_09725_ ), .A2(_05386_ ), .A3(_05462_ ), .A4(_09678_ ), .ZN(_05478_ ) );
OAI21_X1 _20357_ ( .A(\u_lsu.pmem[4355] ), .B1(_03950_ ), .B2(_09468_ ), .ZN(_05479_ ) );
AOI21_X1 _20358_ ( .A(fanout_net_71 ), .B1(_05478_ ), .B2(_05479_ ), .ZN(_02076_ ) );
NAND4_X1 _20359_ ( .A1(_10135_ ), .A2(_05453_ ), .A3(_05427_ ), .A4(_05428_ ), .ZN(_05480_ ) );
OAI21_X1 _20360_ ( .A(\u_lsu.pmem[4034] ), .B1(_10106_ ), .B2(_10110_ ), .ZN(_05481_ ) );
AOI21_X1 _20361_ ( .A(fanout_net_71 ), .B1(_05480_ ), .B2(_05481_ ), .ZN(_02077_ ) );
NAND4_X1 _20362_ ( .A1(_10279_ ), .A2(_05386_ ), .A3(_05462_ ), .A4(_05428_ ), .ZN(_05482_ ) );
OAI21_X1 _20363_ ( .A(\u_lsu.pmem[800] ), .B1(_03335_ ), .B2(_05468_ ), .ZN(_05483_ ) );
AOI21_X1 _20364_ ( .A(fanout_net_71 ), .B1(_05482_ ), .B2(_05483_ ), .ZN(_02078_ ) );
BUF_X4 _20365_ ( .A(_09883_ ), .Z(_05484_ ) );
NAND4_X1 _20366_ ( .A1(_10285_ ), .A2(_05484_ ), .A3(_05462_ ), .A4(_05428_ ), .ZN(_05485_ ) );
OAI21_X1 _20367_ ( .A(\u_lsu.pmem[775] ), .B1(_03347_ ), .B2(_05468_ ), .ZN(_05486_ ) );
AOI21_X1 _20368_ ( .A(fanout_net_71 ), .B1(_05485_ ), .B2(_05486_ ), .ZN(_02079_ ) );
NAND4_X1 _20369_ ( .A1(_10295_ ), .A2(_05484_ ), .A3(_05462_ ), .A4(_05428_ ), .ZN(_05487_ ) );
OAI21_X1 _20370_ ( .A(\u_lsu.pmem[774] ), .B1(_03347_ ), .B2(_05468_ ), .ZN(_05488_ ) );
AOI21_X1 _20371_ ( .A(fanout_net_71 ), .B1(_05487_ ), .B2(_05488_ ), .ZN(_02080_ ) );
NAND4_X1 _20372_ ( .A1(_10299_ ), .A2(_05484_ ), .A3(_05462_ ), .A4(_05428_ ), .ZN(_05489_ ) );
OAI21_X1 _20373_ ( .A(\u_lsu.pmem[773] ), .B1(_03347_ ), .B2(_05468_ ), .ZN(_05490_ ) );
AOI21_X1 _20374_ ( .A(fanout_net_71 ), .B1(_05489_ ), .B2(_05490_ ), .ZN(_02081_ ) );
BUF_X4 _20375_ ( .A(_05166_ ), .Z(_05491_ ) );
NAND4_X1 _20376_ ( .A1(_10306_ ), .A2(_05484_ ), .A3(_05462_ ), .A4(_05491_ ), .ZN(_05492_ ) );
OAI21_X1 _20377_ ( .A(\u_lsu.pmem[772] ), .B1(_03347_ ), .B2(_05468_ ), .ZN(_05493_ ) );
AOI21_X1 _20378_ ( .A(fanout_net_71 ), .B1(_05492_ ), .B2(_05493_ ), .ZN(_02082_ ) );
NAND4_X1 _20379_ ( .A1(_10309_ ), .A2(_05484_ ), .A3(_05462_ ), .A4(_05491_ ), .ZN(_05494_ ) );
OAI21_X1 _20380_ ( .A(\u_lsu.pmem[771] ), .B1(_03347_ ), .B2(_05468_ ), .ZN(_05495_ ) );
AOI21_X1 _20381_ ( .A(fanout_net_71 ), .B1(_05494_ ), .B2(_05495_ ), .ZN(_02083_ ) );
BUF_X4 _20382_ ( .A(_05181_ ), .Z(_05496_ ) );
NAND4_X1 _20383_ ( .A1(_10037_ ), .A2(_05484_ ), .A3(_05496_ ), .A4(_10313_ ), .ZN(_05497_ ) );
BUF_X4 _20384_ ( .A(_09451_ ), .Z(_05498_ ) );
OAI21_X1 _20385_ ( .A(\u_lsu.pmem[770] ), .B1(_03347_ ), .B2(_05498_ ), .ZN(_05499_ ) );
AOI21_X1 _20386_ ( .A(fanout_net_71 ), .B1(_05497_ ), .B2(_05499_ ), .ZN(_02084_ ) );
NAND4_X1 _20387_ ( .A1(_10316_ ), .A2(_05484_ ), .A3(_05496_ ), .A4(_05491_ ), .ZN(_05500_ ) );
OAI21_X1 _20388_ ( .A(\u_lsu.pmem[769] ), .B1(_03347_ ), .B2(_05498_ ), .ZN(_05501_ ) );
AOI21_X1 _20389_ ( .A(fanout_net_71 ), .B1(_05500_ ), .B2(_05501_ ), .ZN(_02085_ ) );
NAND4_X1 _20390_ ( .A1(_10320_ ), .A2(_05484_ ), .A3(_05496_ ), .A4(_05491_ ), .ZN(_05502_ ) );
OAI21_X1 _20391_ ( .A(\u_lsu.pmem[768] ), .B1(_03347_ ), .B2(_05498_ ), .ZN(_05503_ ) );
AOI21_X1 _20392_ ( .A(fanout_net_71 ), .B1(_05502_ ), .B2(_05503_ ), .ZN(_02086_ ) );
NAND4_X1 _20393_ ( .A1(_10037_ ), .A2(_09674_ ), .A3(_04928_ ), .A4(_11245_ ), .ZN(_05504_ ) );
OAI21_X1 _20394_ ( .A(\u_lsu.pmem[743] ), .B1(_03369_ ), .B2(_05498_ ), .ZN(_05505_ ) );
AOI21_X1 _20395_ ( .A(fanout_net_71 ), .B1(_05504_ ), .B2(_05505_ ), .ZN(_02087_ ) );
NAND4_X1 _20396_ ( .A1(_10138_ ), .A2(_05453_ ), .A3(_05427_ ), .A4(_05491_ ), .ZN(_05506_ ) );
OAI21_X1 _20397_ ( .A(\u_lsu.pmem[4033] ), .B1(_10106_ ), .B2(_10110_ ), .ZN(_05507_ ) );
AOI21_X1 _20398_ ( .A(fanout_net_71 ), .B1(_05506_ ), .B2(_05507_ ), .ZN(_02088_ ) );
NAND4_X1 _20399_ ( .A1(_10332_ ), .A2(_05484_ ), .A3(_05496_ ), .A4(_05491_ ), .ZN(_05508_ ) );
OAI21_X1 _20400_ ( .A(\u_lsu.pmem[742] ), .B1(_03369_ ), .B2(_05498_ ), .ZN(_05509_ ) );
AOI21_X1 _20401_ ( .A(fanout_net_71 ), .B1(_05508_ ), .B2(_05509_ ), .ZN(_02089_ ) );
NAND4_X1 _20402_ ( .A1(_10336_ ), .A2(_05484_ ), .A3(_05496_ ), .A4(_05491_ ), .ZN(_05510_ ) );
OAI21_X1 _20403_ ( .A(\u_lsu.pmem[741] ), .B1(_03369_ ), .B2(_05498_ ), .ZN(_05511_ ) );
AOI21_X1 _20404_ ( .A(fanout_net_71 ), .B1(_05510_ ), .B2(_05511_ ), .ZN(_02090_ ) );
BUF_X4 _20405_ ( .A(_09883_ ), .Z(_05512_ ) );
NAND4_X1 _20406_ ( .A1(_10339_ ), .A2(_05512_ ), .A3(_05496_ ), .A4(_05491_ ), .ZN(_05513_ ) );
OAI21_X1 _20407_ ( .A(\u_lsu.pmem[740] ), .B1(_03369_ ), .B2(_05498_ ), .ZN(_05514_ ) );
AOI21_X1 _20408_ ( .A(fanout_net_71 ), .B1(_05513_ ), .B2(_05514_ ), .ZN(_02091_ ) );
NAND4_X1 _20409_ ( .A1(_10345_ ), .A2(_05512_ ), .A3(_05496_ ), .A4(_05491_ ), .ZN(_05515_ ) );
OAI21_X1 _20410_ ( .A(\u_lsu.pmem[739] ), .B1(_03369_ ), .B2(_05498_ ), .ZN(_05516_ ) );
AOI21_X1 _20411_ ( .A(fanout_net_71 ), .B1(_05515_ ), .B2(_05516_ ), .ZN(_02092_ ) );
NAND4_X1 _20412_ ( .A1(_10350_ ), .A2(_05512_ ), .A3(_05496_ ), .A4(_05491_ ), .ZN(_05517_ ) );
OAI21_X1 _20413_ ( .A(\u_lsu.pmem[738] ), .B1(_03369_ ), .B2(_05498_ ), .ZN(_05518_ ) );
AOI21_X1 _20414_ ( .A(fanout_net_71 ), .B1(_05517_ ), .B2(_05518_ ), .ZN(_02093_ ) );
BUF_X4 _20415_ ( .A(_05166_ ), .Z(_05519_ ) );
NAND4_X1 _20416_ ( .A1(_10354_ ), .A2(_05512_ ), .A3(_05496_ ), .A4(_05519_ ), .ZN(_05520_ ) );
OAI21_X1 _20417_ ( .A(\u_lsu.pmem[737] ), .B1(_03369_ ), .B2(_05498_ ), .ZN(_05521_ ) );
AOI21_X1 _20418_ ( .A(fanout_net_72 ), .B1(_05520_ ), .B2(_05521_ ), .ZN(_02094_ ) );
NAND4_X1 _20419_ ( .A1(_10357_ ), .A2(_05512_ ), .A3(_05496_ ), .A4(_05519_ ), .ZN(_05522_ ) );
BUF_X4 _20420_ ( .A(_09451_ ), .Z(_05523_ ) );
OAI21_X1 _20421_ ( .A(\u_lsu.pmem[736] ), .B1(_03369_ ), .B2(_05523_ ), .ZN(_05524_ ) );
AOI21_X1 _20422_ ( .A(fanout_net_72 ), .B1(_05522_ ), .B2(_05524_ ), .ZN(_02095_ ) );
NAND4_X1 _20423_ ( .A1(_10037_ ), .A2(_09674_ ), .A3(_04928_ ), .A4(_11267_ ), .ZN(_05525_ ) );
OAI21_X1 _20424_ ( .A(\u_lsu.pmem[711] ), .B1(_03393_ ), .B2(_05523_ ), .ZN(_05526_ ) );
AOI21_X1 _20425_ ( .A(fanout_net_72 ), .B1(_05525_ ), .B2(_05526_ ), .ZN(_02096_ ) );
BUF_X4 _20426_ ( .A(_05181_ ), .Z(_05527_ ) );
NAND4_X1 _20427_ ( .A1(_10368_ ), .A2(_05512_ ), .A3(_05527_ ), .A4(_05519_ ), .ZN(_05528_ ) );
OAI21_X1 _20428_ ( .A(\u_lsu.pmem[710] ), .B1(_03393_ ), .B2(_05523_ ), .ZN(_05529_ ) );
AOI21_X1 _20429_ ( .A(fanout_net_72 ), .B1(_05528_ ), .B2(_05529_ ), .ZN(_02097_ ) );
NAND4_X1 _20430_ ( .A1(_10371_ ), .A2(_05512_ ), .A3(_05527_ ), .A4(_05519_ ), .ZN(_05530_ ) );
OAI21_X1 _20431_ ( .A(\u_lsu.pmem[709] ), .B1(_03393_ ), .B2(_05523_ ), .ZN(_05531_ ) );
AOI21_X1 _20432_ ( .A(fanout_net_72 ), .B1(_05530_ ), .B2(_05531_ ), .ZN(_02098_ ) );
NAND4_X1 _20433_ ( .A1(_10144_ ), .A2(_05453_ ), .A3(_05427_ ), .A4(_05519_ ), .ZN(_05532_ ) );
OAI21_X1 _20434_ ( .A(\u_lsu.pmem[4032] ), .B1(_10106_ ), .B2(_10110_ ), .ZN(_05533_ ) );
AOI21_X1 _20435_ ( .A(fanout_net_72 ), .B1(_05532_ ), .B2(_05533_ ), .ZN(_02099_ ) );
NAND4_X1 _20436_ ( .A1(_10374_ ), .A2(_05512_ ), .A3(_05527_ ), .A4(_05519_ ), .ZN(_05534_ ) );
OAI21_X1 _20437_ ( .A(\u_lsu.pmem[708] ), .B1(_03393_ ), .B2(_05523_ ), .ZN(_05535_ ) );
AOI21_X1 _20438_ ( .A(fanout_net_72 ), .B1(_05534_ ), .B2(_05535_ ), .ZN(_02100_ ) );
NAND4_X1 _20439_ ( .A1(_10377_ ), .A2(_05512_ ), .A3(_05527_ ), .A4(_05519_ ), .ZN(_05536_ ) );
OAI21_X1 _20440_ ( .A(\u_lsu.pmem[707] ), .B1(_03393_ ), .B2(_05523_ ), .ZN(_05537_ ) );
AOI21_X1 _20441_ ( .A(fanout_net_72 ), .B1(_05536_ ), .B2(_05537_ ), .ZN(_02101_ ) );
NAND4_X1 _20442_ ( .A1(_10381_ ), .A2(_05512_ ), .A3(_05527_ ), .A4(_05519_ ), .ZN(_05538_ ) );
OAI21_X1 _20443_ ( .A(\u_lsu.pmem[706] ), .B1(_03393_ ), .B2(_05523_ ), .ZN(_05539_ ) );
AOI21_X1 _20444_ ( .A(fanout_net_72 ), .B1(_05538_ ), .B2(_05539_ ), .ZN(_02102_ ) );
BUF_X4 _20445_ ( .A(_09883_ ), .Z(_05540_ ) );
NAND4_X1 _20446_ ( .A1(_10384_ ), .A2(_05540_ ), .A3(_05527_ ), .A4(_05519_ ), .ZN(_05541_ ) );
OAI21_X1 _20447_ ( .A(\u_lsu.pmem[705] ), .B1(_03393_ ), .B2(_05523_ ), .ZN(_05542_ ) );
AOI21_X1 _20448_ ( .A(fanout_net_72 ), .B1(_05541_ ), .B2(_05542_ ), .ZN(_02103_ ) );
NAND4_X1 _20449_ ( .A1(_10391_ ), .A2(_05540_ ), .A3(_05527_ ), .A4(_05519_ ), .ZN(_05543_ ) );
OAI21_X1 _20450_ ( .A(\u_lsu.pmem[704] ), .B1(_03393_ ), .B2(_05523_ ), .ZN(_05544_ ) );
AOI21_X1 _20451_ ( .A(fanout_net_72 ), .B1(_05543_ ), .B2(_05544_ ), .ZN(_02104_ ) );
BUF_X4 _20452_ ( .A(_05166_ ), .Z(_05545_ ) );
NAND4_X1 _20453_ ( .A1(_10394_ ), .A2(_05540_ ), .A3(_05527_ ), .A4(_05545_ ), .ZN(_05546_ ) );
OAI21_X1 _20454_ ( .A(\u_lsu.pmem[679] ), .B1(_03417_ ), .B2(_05523_ ), .ZN(_05547_ ) );
AOI21_X1 _20455_ ( .A(fanout_net_72 ), .B1(_05546_ ), .B2(_05547_ ), .ZN(_02105_ ) );
NAND4_X1 _20456_ ( .A1(_10402_ ), .A2(_05540_ ), .A3(_05527_ ), .A4(_05545_ ), .ZN(_05548_ ) );
BUF_X4 _20457_ ( .A(_09451_ ), .Z(_05549_ ) );
OAI21_X1 _20458_ ( .A(\u_lsu.pmem[678] ), .B1(_03417_ ), .B2(_05549_ ), .ZN(_05550_ ) );
AOI21_X1 _20459_ ( .A(fanout_net_72 ), .B1(_05548_ ), .B2(_05550_ ), .ZN(_02106_ ) );
NAND4_X1 _20460_ ( .A1(_10405_ ), .A2(_05540_ ), .A3(_05527_ ), .A4(_05545_ ), .ZN(_05551_ ) );
OAI21_X1 _20461_ ( .A(\u_lsu.pmem[677] ), .B1(_03417_ ), .B2(_05549_ ), .ZN(_05552_ ) );
AOI21_X1 _20462_ ( .A(fanout_net_72 ), .B1(_05551_ ), .B2(_05552_ ), .ZN(_02107_ ) );
BUF_X4 _20463_ ( .A(_05181_ ), .Z(_05553_ ) );
NAND4_X1 _20464_ ( .A1(_10408_ ), .A2(_05540_ ), .A3(_05553_ ), .A4(_05545_ ), .ZN(_05554_ ) );
OAI21_X1 _20465_ ( .A(\u_lsu.pmem[676] ), .B1(_03417_ ), .B2(_05549_ ), .ZN(_05555_ ) );
AOI21_X1 _20466_ ( .A(fanout_net_72 ), .B1(_05554_ ), .B2(_05555_ ), .ZN(_02108_ ) );
NAND4_X1 _20467_ ( .A1(_10411_ ), .A2(_05540_ ), .A3(_05553_ ), .A4(_05545_ ), .ZN(_05556_ ) );
OAI21_X1 _20468_ ( .A(\u_lsu.pmem[675] ), .B1(_03417_ ), .B2(_05549_ ), .ZN(_05557_ ) );
AOI21_X1 _20469_ ( .A(fanout_net_72 ), .B1(_05556_ ), .B2(_05557_ ), .ZN(_02109_ ) );
NAND4_X1 _20470_ ( .A1(_10148_ ), .A2(_05453_ ), .A3(_05427_ ), .A4(_05545_ ), .ZN(_05558_ ) );
INV_X1 _20471_ ( .A(_09494_ ), .ZN(_05559_ ) );
NAND2_X1 _20472_ ( .A1(_05559_ ), .A2(\u_lsu.pmem[4007] ), .ZN(_05560_ ) );
AOI21_X1 _20473_ ( .A(fanout_net_72 ), .B1(_05558_ ), .B2(_05560_ ), .ZN(_02110_ ) );
NAND4_X1 _20474_ ( .A1(_10414_ ), .A2(_05540_ ), .A3(_05553_ ), .A4(_05545_ ), .ZN(_05561_ ) );
OAI21_X1 _20475_ ( .A(\u_lsu.pmem[674] ), .B1(_03417_ ), .B2(_05549_ ), .ZN(_05562_ ) );
AOI21_X1 _20476_ ( .A(fanout_net_72 ), .B1(_05561_ ), .B2(_05562_ ), .ZN(_02111_ ) );
NAND4_X1 _20477_ ( .A1(_10417_ ), .A2(_05540_ ), .A3(_05553_ ), .A4(_05545_ ), .ZN(_05563_ ) );
OAI21_X1 _20478_ ( .A(\u_lsu.pmem[673] ), .B1(_03417_ ), .B2(_05549_ ), .ZN(_05564_ ) );
AOI21_X1 _20479_ ( .A(fanout_net_72 ), .B1(_05563_ ), .B2(_05564_ ), .ZN(_02112_ ) );
NAND4_X1 _20480_ ( .A1(_10037_ ), .A2(_02486_ ), .A3(_03753_ ), .A4(_11292_ ), .ZN(_05565_ ) );
OAI21_X1 _20481_ ( .A(\u_lsu.pmem[672] ), .B1(_03417_ ), .B2(_05549_ ), .ZN(_05566_ ) );
AOI21_X1 _20482_ ( .A(fanout_net_72 ), .B1(_05565_ ), .B2(_05566_ ), .ZN(_02113_ ) );
OAI21_X1 _20483_ ( .A(\u_lsu.pmem[647] ), .B1(_03439_ ), .B2(_05411_ ), .ZN(_05567_ ) );
NAND4_X1 _20484_ ( .A1(_10436_ ), .A2(_04585_ ), .A3(_05401_ ), .A4(_04008_ ), .ZN(_05568_ ) );
AOI21_X1 _20485_ ( .A(fanout_net_72 ), .B1(_05567_ ), .B2(_05568_ ), .ZN(_02114_ ) );
NAND4_X1 _20486_ ( .A1(_03457_ ), .A2(_09658_ ), .A3(_05553_ ), .A4(_05545_ ), .ZN(_05569_ ) );
OAI21_X1 _20487_ ( .A(\u_lsu.pmem[646] ), .B1(_03438_ ), .B2(_05549_ ), .ZN(_05570_ ) );
AOI21_X1 _20488_ ( .A(fanout_net_72 ), .B1(_05569_ ), .B2(_05570_ ), .ZN(_02115_ ) );
NAND4_X1 _20489_ ( .A1(_03457_ ), .A2(_09713_ ), .A3(_03436_ ), .A4(_05545_ ), .ZN(_05571_ ) );
OAI21_X1 _20490_ ( .A(\u_lsu.pmem[645] ), .B1(_03438_ ), .B2(_05549_ ), .ZN(_05572_ ) );
AOI21_X1 _20491_ ( .A(fanout_net_72 ), .B1(_05571_ ), .B2(_05572_ ), .ZN(_02116_ ) );
BUF_X4 _20492_ ( .A(_09515_ ), .Z(_05573_ ) );
NAND4_X1 _20493_ ( .A1(_11320_ ), .A2(_09514_ ), .A3(_05553_ ), .A4(_05573_ ), .ZN(_05574_ ) );
OAI21_X1 _20494_ ( .A(\u_lsu.pmem[644] ), .B1(_03438_ ), .B2(_05549_ ), .ZN(_05575_ ) );
AOI21_X1 _20495_ ( .A(fanout_net_72 ), .B1(_05574_ ), .B2(_05575_ ), .ZN(_02117_ ) );
NAND4_X1 _20496_ ( .A1(_11320_ ), .A2(_09520_ ), .A3(_03436_ ), .A4(_05573_ ), .ZN(_05576_ ) );
BUF_X4 _20497_ ( .A(_09451_ ), .Z(_05577_ ) );
OAI21_X1 _20498_ ( .A(\u_lsu.pmem[643] ), .B1(_03438_ ), .B2(_05577_ ), .ZN(_05578_ ) );
AOI21_X1 _20499_ ( .A(fanout_net_72 ), .B1(_05576_ ), .B2(_05578_ ), .ZN(_02118_ ) );
OAI21_X1 _20500_ ( .A(\u_lsu.pmem[642] ), .B1(_03439_ ), .B2(_05411_ ), .ZN(_05579_ ) );
NAND4_X1 _20501_ ( .A1(_10460_ ), .A2(_04585_ ), .A3(_05401_ ), .A4(_04008_ ), .ZN(_05580_ ) );
AOI21_X1 _20502_ ( .A(fanout_net_72 ), .B1(_05579_ ), .B2(_05580_ ), .ZN(_02119_ ) );
NAND4_X1 _20503_ ( .A1(_11320_ ), .A2(_09544_ ), .A3(_03436_ ), .A4(_05573_ ), .ZN(_05581_ ) );
OAI21_X1 _20504_ ( .A(\u_lsu.pmem[641] ), .B1(_03438_ ), .B2(_05577_ ), .ZN(_05582_ ) );
AOI21_X1 _20505_ ( .A(fanout_net_72 ), .B1(_05581_ ), .B2(_05582_ ), .ZN(_02120_ ) );
NAND4_X1 _20506_ ( .A1(_10156_ ), .A2(_05453_ ), .A3(_05427_ ), .A4(_05573_ ), .ZN(_05583_ ) );
NAND2_X1 _20507_ ( .A1(_05559_ ), .A2(\u_lsu.pmem[4006] ), .ZN(_05584_ ) );
AOI21_X1 _20508_ ( .A(fanout_net_72 ), .B1(_05583_ ), .B2(_05584_ ), .ZN(_02121_ ) );
NAND4_X1 _20509_ ( .A1(_11320_ ), .A2(_09548_ ), .A3(_03436_ ), .A4(_05573_ ), .ZN(_05585_ ) );
OAI21_X1 _20510_ ( .A(\u_lsu.pmem[640] ), .B1(_03438_ ), .B2(_05577_ ), .ZN(_05586_ ) );
AOI21_X1 _20511_ ( .A(fanout_net_72 ), .B1(_05585_ ), .B2(_05586_ ), .ZN(_02122_ ) );
OAI21_X1 _20512_ ( .A(\u_lsu.pmem[615] ), .B1(_03464_ ), .B2(_05411_ ), .ZN(_05587_ ) );
NAND3_X1 _20513_ ( .A1(_09460_ ), .A2(_10330_ ), .A3(_03466_ ), .ZN(_05588_ ) );
AOI21_X1 _20514_ ( .A(fanout_net_72 ), .B1(_05587_ ), .B2(_05588_ ), .ZN(_02123_ ) );
OAI21_X1 _20515_ ( .A(\u_lsu.pmem[614] ), .B1(_03464_ ), .B2(_05411_ ), .ZN(_05589_ ) );
NAND3_X1 _20516_ ( .A1(_09460_ ), .A2(_09579_ ), .A3(_03466_ ), .ZN(_05590_ ) );
AOI21_X1 _20517_ ( .A(fanout_net_73 ), .B1(_05589_ ), .B2(_05590_ ), .ZN(_02124_ ) );
OAI21_X1 _20518_ ( .A(\u_lsu.pmem[613] ), .B1(_03463_ ), .B2(_05411_ ), .ZN(_05591_ ) );
NAND3_X1 _20519_ ( .A1(_09460_ ), .A2(_09586_ ), .A3(_03462_ ), .ZN(_05592_ ) );
AOI21_X1 _20520_ ( .A(fanout_net_73 ), .B1(_05591_ ), .B2(_05592_ ), .ZN(_02125_ ) );
OAI21_X1 _20521_ ( .A(\u_lsu.pmem[612] ), .B1(_03463_ ), .B2(_05411_ ), .ZN(_05593_ ) );
NAND3_X1 _20522_ ( .A1(_09460_ ), .A2(_10486_ ), .A3(_03462_ ), .ZN(_05594_ ) );
AOI21_X1 _20523_ ( .A(fanout_net_73 ), .B1(_05593_ ), .B2(_05594_ ), .ZN(_02126_ ) );
BUF_X4 _20524_ ( .A(_10720_ ), .Z(_05595_ ) );
OAI21_X1 _20525_ ( .A(\u_lsu.pmem[611] ), .B1(_03463_ ), .B2(_05595_ ), .ZN(_05596_ ) );
NAND3_X1 _20526_ ( .A1(_09460_ ), .A2(_09449_ ), .A3(_03462_ ), .ZN(_05597_ ) );
AOI21_X1 _20527_ ( .A(fanout_net_73 ), .B1(_05596_ ), .B2(_05597_ ), .ZN(_02127_ ) );
OAI21_X1 _20528_ ( .A(\u_lsu.pmem[610] ), .B1(_03463_ ), .B2(_05595_ ), .ZN(_05598_ ) );
NAND3_X1 _20529_ ( .A1(_09460_ ), .A2(_09695_ ), .A3(_03462_ ), .ZN(_05599_ ) );
AOI21_X1 _20530_ ( .A(fanout_net_73 ), .B1(_05598_ ), .B2(_05599_ ), .ZN(_02128_ ) );
OAI21_X1 _20531_ ( .A(\u_lsu.pmem[609] ), .B1(_03463_ ), .B2(_05595_ ), .ZN(_05600_ ) );
NAND3_X1 _20532_ ( .A1(_09460_ ), .A2(_09698_ ), .A3(_03462_ ), .ZN(_05601_ ) );
AOI21_X1 _20533_ ( .A(fanout_net_73 ), .B1(_05600_ ), .B2(_05601_ ), .ZN(_02129_ ) );
OAI21_X1 _20534_ ( .A(\u_lsu.pmem[608] ), .B1(_03463_ ), .B2(_05595_ ), .ZN(_05602_ ) );
NAND3_X1 _20535_ ( .A1(_09460_ ), .A2(_09622_ ), .A3(_03462_ ), .ZN(_05603_ ) );
AOI21_X1 _20536_ ( .A(fanout_net_73 ), .B1(_05602_ ), .B2(_05603_ ), .ZN(_02130_ ) );
OAI21_X1 _20537_ ( .A(\u_lsu.pmem[583] ), .B1(_03488_ ), .B2(_05595_ ), .ZN(_05604_ ) );
NAND4_X1 _20538_ ( .A1(_03957_ ), .A2(_09477_ ), .A3(_09741_ ), .A4(_03499_ ), .ZN(_05605_ ) );
AOI21_X1 _20539_ ( .A(fanout_net_73 ), .B1(_05604_ ), .B2(_05605_ ), .ZN(_02131_ ) );
NAND4_X1 _20540_ ( .A1(_10160_ ), .A2(_05453_ ), .A3(_05427_ ), .A4(_05573_ ), .ZN(_05606_ ) );
NAND2_X1 _20541_ ( .A1(_05559_ ), .A2(\u_lsu.pmem[4005] ), .ZN(_05607_ ) );
AOI21_X1 _20542_ ( .A(fanout_net_73 ), .B1(_05606_ ), .B2(_05607_ ), .ZN(_02132_ ) );
OAI21_X1 _20543_ ( .A(\u_lsu.pmem[582] ), .B1(_03488_ ), .B2(_05595_ ), .ZN(_05608_ ) );
NAND4_X1 _20544_ ( .A1(_03957_ ), .A2(_09477_ ), .A3(_09578_ ), .A4(_03499_ ), .ZN(_05609_ ) );
AOI21_X1 _20545_ ( .A(fanout_net_73 ), .B1(_05608_ ), .B2(_05609_ ), .ZN(_02133_ ) );
OAI21_X1 _20546_ ( .A(\u_lsu.pmem[581] ), .B1(_03487_ ), .B2(_05595_ ), .ZN(_05610_ ) );
NAND4_X1 _20547_ ( .A1(_09444_ ), .A2(_09477_ ), .A3(_09585_ ), .A4(_03499_ ), .ZN(_05611_ ) );
AOI21_X1 _20548_ ( .A(fanout_net_73 ), .B1(_05610_ ), .B2(_05611_ ), .ZN(_02134_ ) );
OAI21_X1 _20549_ ( .A(\u_lsu.pmem[580] ), .B1(_03487_ ), .B2(_05595_ ), .ZN(_05612_ ) );
NAND4_X1 _20550_ ( .A1(_09444_ ), .A2(_09477_ ), .A3(_11151_ ), .A4(_03499_ ), .ZN(_05613_ ) );
AOI21_X1 _20551_ ( .A(fanout_net_73 ), .B1(_05612_ ), .B2(_05613_ ), .ZN(_02135_ ) );
OAI21_X1 _20552_ ( .A(\u_lsu.pmem[579] ), .B1(_03487_ ), .B2(_05595_ ), .ZN(_05614_ ) );
NAND4_X1 _20553_ ( .A1(_09444_ ), .A2(_09477_ ), .A3(_09448_ ), .A4(_03499_ ), .ZN(_05615_ ) );
AOI21_X1 _20554_ ( .A(fanout_net_73 ), .B1(_05614_ ), .B2(_05615_ ), .ZN(_02136_ ) );
OAI21_X1 _20555_ ( .A(\u_lsu.pmem[578] ), .B1(_03487_ ), .B2(_05595_ ), .ZN(_05616_ ) );
NAND4_X1 _20556_ ( .A1(_09444_ ), .A2(_09477_ ), .A3(_10015_ ), .A4(_03499_ ), .ZN(_05617_ ) );
AOI21_X1 _20557_ ( .A(fanout_net_73 ), .B1(_05616_ ), .B2(_05617_ ), .ZN(_02137_ ) );
BUF_X4 _20558_ ( .A(_10720_ ), .Z(_05618_ ) );
OAI21_X1 _20559_ ( .A(\u_lsu.pmem[577] ), .B1(_03487_ ), .B2(_05618_ ), .ZN(_05619_ ) );
NAND4_X1 _20560_ ( .A1(_09444_ ), .A2(_09477_ ), .A3(_09616_ ), .A4(_11369_ ), .ZN(_05620_ ) );
AOI21_X1 _20561_ ( .A(fanout_net_73 ), .B1(_05619_ ), .B2(_05620_ ), .ZN(_02138_ ) );
OAI21_X1 _20562_ ( .A(\u_lsu.pmem[576] ), .B1(_03487_ ), .B2(_05618_ ), .ZN(_05621_ ) );
NAND4_X1 _20563_ ( .A1(_09444_ ), .A2(_09477_ ), .A3(_09621_ ), .A4(_11369_ ), .ZN(_05622_ ) );
AOI21_X1 _20564_ ( .A(fanout_net_73 ), .B1(_05621_ ), .B2(_05622_ ), .ZN(_02139_ ) );
NAND4_X1 _20565_ ( .A1(_10527_ ), .A2(_05540_ ), .A3(_05553_ ), .A4(_05573_ ), .ZN(_05623_ ) );
OAI21_X1 _20566_ ( .A(\u_lsu.pmem[551] ), .B1(_03519_ ), .B2(_05577_ ), .ZN(_05624_ ) );
AOI21_X1 _20567_ ( .A(fanout_net_73 ), .B1(_05623_ ), .B2(_05624_ ), .ZN(_02140_ ) );
BUF_X4 _20568_ ( .A(_09883_ ), .Z(_05625_ ) );
NAND4_X1 _20569_ ( .A1(_10535_ ), .A2(_05625_ ), .A3(_05553_ ), .A4(_05573_ ), .ZN(_05626_ ) );
OAI21_X1 _20570_ ( .A(\u_lsu.pmem[550] ), .B1(_03519_ ), .B2(_05577_ ), .ZN(_05627_ ) );
AOI21_X1 _20571_ ( .A(fanout_net_73 ), .B1(_05626_ ), .B2(_05627_ ), .ZN(_02141_ ) );
NAND4_X1 _20572_ ( .A1(_10538_ ), .A2(_05625_ ), .A3(_05553_ ), .A4(_05573_ ), .ZN(_05628_ ) );
OAI21_X1 _20573_ ( .A(\u_lsu.pmem[549] ), .B1(_03519_ ), .B2(_05577_ ), .ZN(_05629_ ) );
AOI21_X1 _20574_ ( .A(fanout_net_73 ), .B1(_05628_ ), .B2(_05629_ ), .ZN(_02142_ ) );
NAND4_X1 _20575_ ( .A1(_10166_ ), .A2(_05453_ ), .A3(_05427_ ), .A4(_05573_ ), .ZN(_05630_ ) );
NAND2_X1 _20576_ ( .A1(_05559_ ), .A2(\u_lsu.pmem[4004] ), .ZN(_05631_ ) );
AOI21_X1 _20577_ ( .A(fanout_net_73 ), .B1(_05630_ ), .B2(_05631_ ), .ZN(_02143_ ) );
NAND3_X1 _20578_ ( .A1(_05448_ ), .A2(_11152_ ), .A3(_03512_ ), .ZN(_05632_ ) );
OAI21_X1 _20579_ ( .A(\u_lsu.pmem[548] ), .B1(_03519_ ), .B2(_05577_ ), .ZN(_05633_ ) );
AOI21_X1 _20580_ ( .A(fanout_net_73 ), .B1(_05632_ ), .B2(_05633_ ), .ZN(_02144_ ) );
NAND3_X1 _20581_ ( .A1(_05448_ ), .A2(_11155_ ), .A3(_03512_ ), .ZN(_05634_ ) );
OAI21_X1 _20582_ ( .A(\u_lsu.pmem[547] ), .B1(_03519_ ), .B2(_05577_ ), .ZN(_05635_ ) );
AOI21_X1 _20583_ ( .A(fanout_net_73 ), .B1(_05634_ ), .B2(_05635_ ), .ZN(_02145_ ) );
NAND3_X1 _20584_ ( .A1(_09573_ ), .A2(_11158_ ), .A3(_03512_ ), .ZN(_05636_ ) );
OAI21_X1 _20585_ ( .A(\u_lsu.pmem[546] ), .B1(_03519_ ), .B2(_05577_ ), .ZN(_05637_ ) );
AOI21_X1 _20586_ ( .A(fanout_net_73 ), .B1(_05636_ ), .B2(_05637_ ), .ZN(_02146_ ) );
NAND3_X1 _20587_ ( .A1(_09573_ ), .A2(_11163_ ), .A3(_03512_ ), .ZN(_05638_ ) );
OAI21_X1 _20588_ ( .A(\u_lsu.pmem[545] ), .B1(_03519_ ), .B2(_05577_ ), .ZN(_05639_ ) );
AOI21_X1 _20589_ ( .A(fanout_net_73 ), .B1(_05638_ ), .B2(_05639_ ), .ZN(_02147_ ) );
BUF_X4 _20590_ ( .A(_09515_ ), .Z(_05640_ ) );
NAND4_X1 _20591_ ( .A1(_10556_ ), .A2(_05625_ ), .A3(_05553_ ), .A4(_05640_ ), .ZN(_05641_ ) );
BUF_X4 _20592_ ( .A(_09451_ ), .Z(_05642_ ) );
OAI21_X1 _20593_ ( .A(\u_lsu.pmem[544] ), .B1(_03519_ ), .B2(_05642_ ), .ZN(_05643_ ) );
AOI21_X1 _20594_ ( .A(fanout_net_73 ), .B1(_05641_ ), .B2(_05643_ ), .ZN(_02148_ ) );
OAI21_X1 _20595_ ( .A(\u_lsu.pmem[519] ), .B1(_03532_ ), .B2(_05618_ ), .ZN(_05644_ ) );
NAND3_X1 _20596_ ( .A1(_03534_ ), .A2(_11423_ ), .A3(_03950_ ), .ZN(_05645_ ) );
AOI21_X1 _20597_ ( .A(fanout_net_73 ), .B1(_05644_ ), .B2(_05645_ ), .ZN(_02149_ ) );
OAI21_X1 _20598_ ( .A(\u_lsu.pmem[518] ), .B1(_03532_ ), .B2(_05618_ ), .ZN(_05646_ ) );
NAND3_X1 _20599_ ( .A1(_03534_ ), .A2(_10444_ ), .A3(_03950_ ), .ZN(_05647_ ) );
AOI21_X1 _20600_ ( .A(fanout_net_73 ), .B1(_05646_ ), .B2(_05647_ ), .ZN(_02150_ ) );
OAI21_X1 _20601_ ( .A(\u_lsu.pmem[517] ), .B1(_03532_ ), .B2(_05618_ ), .ZN(_05648_ ) );
NAND3_X1 _20602_ ( .A1(_03534_ ), .A2(_10448_ ), .A3(_03950_ ), .ZN(_05649_ ) );
AOI21_X1 _20603_ ( .A(fanout_net_73 ), .B1(_05648_ ), .B2(_05649_ ), .ZN(_02151_ ) );
OAI21_X1 _20604_ ( .A(\u_lsu.pmem[516] ), .B1(_03532_ ), .B2(_05618_ ), .ZN(_05650_ ) );
NAND3_X1 _20605_ ( .A1(_03534_ ), .A2(_10453_ ), .A3(_03950_ ), .ZN(_05651_ ) );
AOI21_X1 _20606_ ( .A(fanout_net_73 ), .B1(_05650_ ), .B2(_05651_ ), .ZN(_02152_ ) );
NAND4_X1 _20607_ ( .A1(_10575_ ), .A2(_09676_ ), .A3(_09540_ ), .A4(_05011_ ), .ZN(_05652_ ) );
OAI21_X1 _20608_ ( .A(\u_lsu.pmem[515] ), .B1(_03531_ ), .B2(_05642_ ), .ZN(_05653_ ) );
AOI21_X1 _20609_ ( .A(fanout_net_73 ), .B1(_05652_ ), .B2(_05653_ ), .ZN(_02153_ ) );
NAND4_X1 _20610_ ( .A1(_10169_ ), .A2(_05453_ ), .A3(_05427_ ), .A4(_05640_ ), .ZN(_05654_ ) );
NAND2_X1 _20611_ ( .A1(_05559_ ), .A2(\u_lsu.pmem[4003] ), .ZN(_05655_ ) );
AOI21_X1 _20612_ ( .A(fanout_net_74 ), .B1(_05654_ ), .B2(_05655_ ), .ZN(_02154_ ) );
BUF_X4 _20613_ ( .A(_09476_ ), .Z(_05656_ ) );
NAND4_X1 _20614_ ( .A1(_10584_ ), .A2(_09806_ ), .A3(_05656_ ), .A4(_05640_ ), .ZN(_05657_ ) );
OAI21_X1 _20615_ ( .A(\u_lsu.pmem[514] ), .B1(_03531_ ), .B2(_05642_ ), .ZN(_05658_ ) );
AOI21_X1 _20616_ ( .A(fanout_net_74 ), .B1(_05657_ ), .B2(_05658_ ), .ZN(_02155_ ) );
OAI21_X1 _20617_ ( .A(\u_lsu.pmem[513] ), .B1(_03532_ ), .B2(_05618_ ), .ZN(_05659_ ) );
NAND3_X1 _20618_ ( .A1(_03534_ ), .A2(_10463_ ), .A3(_03950_ ), .ZN(_05660_ ) );
AOI21_X1 _20619_ ( .A(fanout_net_74 ), .B1(_05659_ ), .B2(_05660_ ), .ZN(_02156_ ) );
NAND4_X1 _20620_ ( .A1(_10591_ ), .A2(_09676_ ), .A3(_09540_ ), .A4(_05011_ ), .ZN(_05661_ ) );
OAI21_X1 _20621_ ( .A(\u_lsu.pmem[512] ), .B1(_03531_ ), .B2(_05642_ ), .ZN(_05662_ ) );
AOI21_X1 _20622_ ( .A(fanout_net_74 ), .B1(_05661_ ), .B2(_05662_ ), .ZN(_02157_ ) );
NAND4_X1 _20623_ ( .A1(_10037_ ), .A2(_09674_ ), .A3(_09741_ ), .A4(_11442_ ), .ZN(_05663_ ) );
OAI21_X1 _20624_ ( .A(\u_lsu.pmem[487] ), .B1(_03556_ ), .B2(_05642_ ), .ZN(_05664_ ) );
AOI21_X1 _20625_ ( .A(fanout_net_74 ), .B1(_05663_ ), .B2(_05664_ ), .ZN(_02158_ ) );
NAND4_X1 _20626_ ( .A1(_10603_ ), .A2(_05625_ ), .A3(_05656_ ), .A4(_05640_ ), .ZN(_05665_ ) );
OAI21_X1 _20627_ ( .A(\u_lsu.pmem[486] ), .B1(_03556_ ), .B2(_05642_ ), .ZN(_05666_ ) );
AOI21_X1 _20628_ ( .A(fanout_net_74 ), .B1(_05665_ ), .B2(_05666_ ), .ZN(_02159_ ) );
NAND4_X1 _20629_ ( .A1(_10608_ ), .A2(_05625_ ), .A3(_05656_ ), .A4(_05640_ ), .ZN(_05667_ ) );
OAI21_X1 _20630_ ( .A(\u_lsu.pmem[485] ), .B1(_03556_ ), .B2(_05642_ ), .ZN(_05668_ ) );
AOI21_X1 _20631_ ( .A(fanout_net_74 ), .B1(_05667_ ), .B2(_05668_ ), .ZN(_02160_ ) );
NAND4_X1 _20632_ ( .A1(_10611_ ), .A2(_05625_ ), .A3(_05656_ ), .A4(_05640_ ), .ZN(_05669_ ) );
OAI21_X1 _20633_ ( .A(\u_lsu.pmem[484] ), .B1(_03556_ ), .B2(_05642_ ), .ZN(_05670_ ) );
AOI21_X1 _20634_ ( .A(fanout_net_74 ), .B1(_05669_ ), .B2(_05670_ ), .ZN(_02161_ ) );
NAND4_X1 _20635_ ( .A1(_10614_ ), .A2(_05625_ ), .A3(_05656_ ), .A4(_05640_ ), .ZN(_05671_ ) );
OAI21_X1 _20636_ ( .A(\u_lsu.pmem[483] ), .B1(_03556_ ), .B2(_05642_ ), .ZN(_05672_ ) );
AOI21_X1 _20637_ ( .A(fanout_net_74 ), .B1(_05671_ ), .B2(_05672_ ), .ZN(_02162_ ) );
NAND4_X1 _20638_ ( .A1(_10617_ ), .A2(_05625_ ), .A3(_05656_ ), .A4(_05640_ ), .ZN(_05673_ ) );
OAI21_X1 _20639_ ( .A(\u_lsu.pmem[482] ), .B1(_03556_ ), .B2(_05642_ ), .ZN(_05674_ ) );
AOI21_X1 _20640_ ( .A(fanout_net_74 ), .B1(_05673_ ), .B2(_05674_ ), .ZN(_02163_ ) );
NAND4_X1 _20641_ ( .A1(_10621_ ), .A2(_05625_ ), .A3(_05656_ ), .A4(_05640_ ), .ZN(_05675_ ) );
BUF_X4 _20642_ ( .A(_09451_ ), .Z(_05676_ ) );
OAI21_X1 _20643_ ( .A(\u_lsu.pmem[481] ), .B1(_03556_ ), .B2(_05676_ ), .ZN(_05677_ ) );
AOI21_X1 _20644_ ( .A(fanout_net_74 ), .B1(_05675_ ), .B2(_05677_ ), .ZN(_02164_ ) );
NAND4_X1 _20645_ ( .A1(_10172_ ), .A2(_05453_ ), .A3(_10579_ ), .A4(_05640_ ), .ZN(_05678_ ) );
NAND2_X1 _20646_ ( .A1(_05559_ ), .A2(\u_lsu.pmem[4002] ), .ZN(_05679_ ) );
AOI21_X1 _20647_ ( .A(fanout_net_74 ), .B1(_05678_ ), .B2(_05679_ ), .ZN(_02165_ ) );
BUF_X4 _20648_ ( .A(_09515_ ), .Z(_05680_ ) );
NAND4_X1 _20649_ ( .A1(_10624_ ), .A2(_05625_ ), .A3(_05656_ ), .A4(_05680_ ), .ZN(_05681_ ) );
OAI21_X1 _20650_ ( .A(\u_lsu.pmem[480] ), .B1(_03556_ ), .B2(_05676_ ), .ZN(_05682_ ) );
AOI21_X1 _20651_ ( .A(fanout_net_74 ), .B1(_05681_ ), .B2(_05682_ ), .ZN(_02166_ ) );
NAND4_X1 _20652_ ( .A1(_10037_ ), .A2(_09674_ ), .A3(_09741_ ), .A4(_11469_ ), .ZN(_05683_ ) );
OAI21_X1 _20653_ ( .A(\u_lsu.pmem[455] ), .B1(_03583_ ), .B2(_05676_ ), .ZN(_05684_ ) );
AOI21_X1 _20654_ ( .A(fanout_net_74 ), .B1(_05683_ ), .B2(_05684_ ), .ZN(_02167_ ) );
BUF_X4 _20655_ ( .A(_09883_ ), .Z(_05685_ ) );
NAND4_X1 _20656_ ( .A1(_10632_ ), .A2(_05685_ ), .A3(_05656_ ), .A4(_05680_ ), .ZN(_05686_ ) );
OAI21_X1 _20657_ ( .A(\u_lsu.pmem[454] ), .B1(_03583_ ), .B2(_05676_ ), .ZN(_05687_ ) );
AOI21_X1 _20658_ ( .A(fanout_net_74 ), .B1(_05686_ ), .B2(_05687_ ), .ZN(_02168_ ) );
NAND4_X1 _20659_ ( .A1(_10635_ ), .A2(_05685_ ), .A3(_05656_ ), .A4(_05680_ ), .ZN(_05688_ ) );
OAI21_X1 _20660_ ( .A(\u_lsu.pmem[453] ), .B1(_03583_ ), .B2(_05676_ ), .ZN(_05689_ ) );
AOI21_X1 _20661_ ( .A(fanout_net_74 ), .B1(_05688_ ), .B2(_05689_ ), .ZN(_02169_ ) );
BUF_X4 _20662_ ( .A(_09476_ ), .Z(_05690_ ) );
NAND4_X1 _20663_ ( .A1(_10641_ ), .A2(_05685_ ), .A3(_05690_ ), .A4(_05680_ ), .ZN(_05691_ ) );
OAI21_X1 _20664_ ( .A(\u_lsu.pmem[452] ), .B1(_03583_ ), .B2(_05676_ ), .ZN(_05692_ ) );
AOI21_X1 _20665_ ( .A(fanout_net_74 ), .B1(_05691_ ), .B2(_05692_ ), .ZN(_02170_ ) );
NAND4_X1 _20666_ ( .A1(_10645_ ), .A2(_05685_ ), .A3(_05690_ ), .A4(_05680_ ), .ZN(_05693_ ) );
OAI21_X1 _20667_ ( .A(\u_lsu.pmem[451] ), .B1(_03583_ ), .B2(_05676_ ), .ZN(_05694_ ) );
AOI21_X1 _20668_ ( .A(fanout_net_74 ), .B1(_05693_ ), .B2(_05694_ ), .ZN(_02171_ ) );
NAND4_X1 _20669_ ( .A1(_10649_ ), .A2(_05685_ ), .A3(_05690_ ), .A4(_05680_ ), .ZN(_05695_ ) );
OAI21_X1 _20670_ ( .A(\u_lsu.pmem[450] ), .B1(_03583_ ), .B2(_05676_ ), .ZN(_05696_ ) );
AOI21_X1 _20671_ ( .A(fanout_net_74 ), .B1(_05695_ ), .B2(_05696_ ), .ZN(_02172_ ) );
NAND4_X1 _20672_ ( .A1(_10652_ ), .A2(_05685_ ), .A3(_05690_ ), .A4(_05680_ ), .ZN(_05697_ ) );
OAI21_X1 _20673_ ( .A(\u_lsu.pmem[449] ), .B1(_03583_ ), .B2(_05676_ ), .ZN(_05698_ ) );
AOI21_X1 _20674_ ( .A(fanout_net_74 ), .B1(_05697_ ), .B2(_05698_ ), .ZN(_02173_ ) );
NAND4_X1 _20675_ ( .A1(_10655_ ), .A2(_05685_ ), .A3(_05690_ ), .A4(_05680_ ), .ZN(_05699_ ) );
OAI21_X1 _20676_ ( .A(\u_lsu.pmem[448] ), .B1(_03583_ ), .B2(_05676_ ), .ZN(_05700_ ) );
AOI21_X1 _20677_ ( .A(fanout_net_74 ), .B1(_05699_ ), .B2(_05700_ ), .ZN(_02174_ ) );
NAND4_X1 _20678_ ( .A1(_10658_ ), .A2(_05685_ ), .A3(_05690_ ), .A4(_05680_ ), .ZN(_05701_ ) );
OAI21_X1 _20679_ ( .A(\u_lsu.pmem[423] ), .B1(_03608_ ), .B2(_09452_ ), .ZN(_05702_ ) );
AOI21_X1 _20680_ ( .A(fanout_net_74 ), .B1(_05701_ ), .B2(_05702_ ), .ZN(_02175_ ) );
NAND4_X1 _20681_ ( .A1(_10176_ ), .A2(_03673_ ), .A3(_10579_ ), .A4(_05680_ ), .ZN(_05703_ ) );
NAND2_X1 _20682_ ( .A1(_05559_ ), .A2(\u_lsu.pmem[4001] ), .ZN(_05704_ ) );
AOI21_X1 _20683_ ( .A(fanout_net_74 ), .B1(_05703_ ), .B2(_05704_ ), .ZN(_02176_ ) );
NAND4_X1 _20684_ ( .A1(_10665_ ), .A2(_05685_ ), .A3(_05690_ ), .A4(_10446_ ), .ZN(_05705_ ) );
OAI21_X1 _20685_ ( .A(\u_lsu.pmem[422] ), .B1(_03608_ ), .B2(_09452_ ), .ZN(_05706_ ) );
AOI21_X1 _20686_ ( .A(fanout_net_74 ), .B1(_05705_ ), .B2(_05706_ ), .ZN(_02177_ ) );
NAND4_X1 _20687_ ( .A1(_10668_ ), .A2(_05685_ ), .A3(_05690_ ), .A4(_10446_ ), .ZN(_05707_ ) );
OAI21_X1 _20688_ ( .A(\u_lsu.pmem[421] ), .B1(_03608_ ), .B2(_09452_ ), .ZN(_05708_ ) );
AOI21_X1 _20689_ ( .A(fanout_net_74 ), .B1(_05707_ ), .B2(_05708_ ), .ZN(_02178_ ) );
NAND4_X1 _20690_ ( .A1(_10671_ ), .A2(_09884_ ), .A3(_05690_ ), .A4(_10446_ ), .ZN(_05709_ ) );
OAI21_X1 _20691_ ( .A(\u_lsu.pmem[420] ), .B1(_03608_ ), .B2(_09452_ ), .ZN(_05710_ ) );
AOI21_X1 _20692_ ( .A(fanout_net_74 ), .B1(_05709_ ), .B2(_05710_ ), .ZN(_02179_ ) );
NAND4_X1 _20693_ ( .A1(_10674_ ), .A2(_09884_ ), .A3(_05690_ ), .A4(_10446_ ), .ZN(_05711_ ) );
OAI21_X1 _20694_ ( .A(\u_lsu.pmem[419] ), .B1(_03608_ ), .B2(_09452_ ), .ZN(_05712_ ) );
AOI21_X1 _20695_ ( .A(fanout_net_74 ), .B1(_05711_ ), .B2(_05712_ ), .ZN(_02180_ ) );
NAND4_X1 _20696_ ( .A1(_10679_ ), .A2(_09884_ ), .A3(_09885_ ), .A4(_10446_ ), .ZN(_05713_ ) );
OAI21_X1 _20697_ ( .A(\u_lsu.pmem[418] ), .B1(_03608_ ), .B2(_09452_ ), .ZN(_05714_ ) );
AOI21_X1 _20698_ ( .A(fanout_net_74 ), .B1(_05713_ ), .B2(_05714_ ), .ZN(_02181_ ) );
NAND4_X1 _20699_ ( .A1(_10682_ ), .A2(_09884_ ), .A3(_09885_ ), .A4(_10446_ ), .ZN(_05715_ ) );
OAI21_X1 _20700_ ( .A(\u_lsu.pmem[417] ), .B1(_03608_ ), .B2(_09452_ ), .ZN(_05716_ ) );
AOI21_X1 _20701_ ( .A(fanout_net_74 ), .B1(_05715_ ), .B2(_05716_ ), .ZN(_02182_ ) );
NAND4_X1 _20702_ ( .A1(_10037_ ), .A2(_09674_ ), .A3(_09621_ ), .A4(_11499_ ), .ZN(_05717_ ) );
OAI21_X1 _20703_ ( .A(\u_lsu.pmem[416] ), .B1(_03608_ ), .B2(_09452_ ), .ZN(_05718_ ) );
AOI21_X1 _20704_ ( .A(fanout_net_74 ), .B1(_05717_ ), .B2(_05718_ ), .ZN(_02183_ ) );
OAI21_X1 _20705_ ( .A(\u_lsu.pmem[391] ), .B1(_09508_ ), .B2(_05618_ ), .ZN(_05719_ ) );
NAND4_X1 _20706_ ( .A1(_09512_ ), .A2(_08582_ ), .A3(_09456_ ), .A4(_04008_ ), .ZN(_05720_ ) );
AOI21_X1 _20707_ ( .A(fanout_net_75 ), .B1(_05719_ ), .B2(_05720_ ), .ZN(_02184_ ) );
OAI21_X1 _20708_ ( .A(\u_lsu.pmem[390] ), .B1(_09508_ ), .B2(_05618_ ), .ZN(_05721_ ) );
NAND4_X1 _20709_ ( .A1(_09512_ ), .A2(_09575_ ), .A3(_09456_ ), .A4(_04008_ ), .ZN(_05722_ ) );
AOI21_X1 _20710_ ( .A(fanout_net_75 ), .B1(_05721_ ), .B2(_05722_ ), .ZN(_02185_ ) );
OAI21_X1 _20711_ ( .A(\u_lsu.pmem[389] ), .B1(_09508_ ), .B2(_05618_ ), .ZN(_05723_ ) );
NAND4_X1 _20712_ ( .A1(_09512_ ), .A2(_09582_ ), .A3(_09456_ ), .A4(_04008_ ), .ZN(_05724_ ) );
AOI21_X1 _20713_ ( .A(fanout_net_75 ), .B1(_05723_ ), .B2(_05724_ ), .ZN(_02186_ ) );
NAND2_X1 _20714_ ( .A1(_09429_ ), .A2(_08908_ ), .ZN(_05725_ ) );
AND2_X1 _20715_ ( .A1(_08944_ ), .A2(_08997_ ), .ZN(_05726_ ) );
INV_X1 _20716_ ( .A(_05726_ ), .ZN(_05727_ ) );
OAI21_X1 _20717_ ( .A(_08902_ ), .B1(\ifu_rdata[4] ), .B2(_08903_ ), .ZN(_05728_ ) );
NOR2_X1 _20718_ ( .A1(_05727_ ), .A2(_05728_ ), .ZN(_05729_ ) );
INV_X1 _20719_ ( .A(_05729_ ), .ZN(_05730_ ) );
BUF_X4 _20720_ ( .A(_05730_ ), .Z(_05731_ ) );
OAI21_X1 _20721_ ( .A(_05725_ ), .B1(_09439_ ), .B2(_05731_ ), .ZN(_05732_ ) );
NOR3_X1 _20722_ ( .A1(\ifu_rdata[2] ), .A2(\ifu_rdata[4] ), .A3(\ifu_rdata[5] ), .ZN(_05733_ ) );
AND2_X2 _20723_ ( .A1(_05733_ ), .A2(_08902_ ), .ZN(_05734_ ) );
INV_X1 _20724_ ( .A(_05734_ ), .ZN(_05735_ ) );
OAI21_X1 _20725_ ( .A(_05735_ ), .B1(_09439_ ), .B2(_08913_ ), .ZN(_05736_ ) );
INV_X1 _20726_ ( .A(_09081_ ), .ZN(_05737_ ) );
AND3_X1 _20727_ ( .A1(_10428_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_09089_ ), .ZN(_05738_ ) );
BUF_X4 _20728_ ( .A(_09111_ ), .Z(_05739_ ) );
BUF_X4 _20729_ ( .A(_09551_ ), .Z(_05740_ ) );
AOI221_X2 _20730_ ( .A(_05738_ ), .B1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_05739_ ), .C1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_05740_ ), .ZN(_05741_ ) );
NAND3_X1 _20731_ ( .A1(_09067_ ), .A2(_09091_ ), .A3(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05742_ ) );
AOI21_X1 _20732_ ( .A(_05737_ ), .B1(_05741_ ), .B2(_05742_ ), .ZN(_05743_ ) );
BUF_X4 _20733_ ( .A(_05737_ ), .Z(_05744_ ) );
BUF_X4 _20734_ ( .A(_09089_ ), .Z(_05745_ ) );
MUX2_X1 _20735_ ( .A(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .S(_05745_ ), .Z(_05746_ ) );
MUX2_X1 _20736_ ( .A(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .S(_05745_ ), .Z(_05747_ ) );
BUF_X2 _20737_ ( .A(_10428_ ), .Z(_05748_ ) );
MUX2_X1 _20738_ ( .A(_05746_ ), .B(_05747_ ), .S(_05748_ ), .Z(_05749_ ) );
AOI211_X1 _20739_ ( .A(_09053_ ), .B(_05743_ ), .C1(_05744_ ), .C2(_05749_ ), .ZN(_05750_ ) );
BUF_X4 _20740_ ( .A(_05737_ ), .Z(_05751_ ) );
BUF_X4 _20741_ ( .A(_09625_ ), .Z(_05752_ ) );
AOI22_X1 _20742_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_09552_ ), .B1(_05752_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05753_ ) );
AOI22_X1 _20743_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_09121_ ), .B1(_09526_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05754_ ) );
AOI21_X1 _20744_ ( .A(_05751_ ), .B1(_05753_ ), .B2(_05754_ ), .ZN(_05755_ ) );
AOI22_X1 _20745_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_09552_ ), .B1(_05752_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05756_ ) );
AOI22_X1 _20746_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_09121_ ), .B1(_09526_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05757_ ) );
AOI21_X1 _20747_ ( .A(_09082_ ), .B1(_05756_ ), .B2(_05757_ ), .ZN(_05758_ ) );
NOR3_X1 _20748_ ( .A1(_09479_ ), .A2(_05755_ ), .A3(_05758_ ), .ZN(_05759_ ) );
NOR3_X1 _20749_ ( .A1(_05750_ ), .A2(_09045_ ), .A3(_05759_ ), .ZN(_05760_ ) );
BUF_X4 _20750_ ( .A(_09625_ ), .Z(_05761_ ) );
BUF_X4 _20751_ ( .A(_09121_ ), .Z(_05762_ ) );
AOI22_X1 _20752_ ( .A1(_05761_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_05762_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_05763_ ) );
BUF_X4 _20753_ ( .A(_09067_ ), .Z(_05764_ ) );
BUF_X4 _20754_ ( .A(_05745_ ), .Z(_05765_ ) );
BUF_X4 _20755_ ( .A(_05765_ ), .Z(_05766_ ) );
NAND3_X1 _20756_ ( .A1(_05764_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_05766_ ), .ZN(_05767_ ) );
BUF_X4 _20757_ ( .A(_08970_ ), .Z(_05768_ ) );
BUF_X4 _20758_ ( .A(_09065_ ), .Z(_05769_ ) );
OAI211_X1 _20759_ ( .A(_09091_ ), .B(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_05768_ ), .C2(_05769_ ), .ZN(_05770_ ) );
NAND4_X1 _20760_ ( .A1(_05763_ ), .A2(_05751_ ), .A3(_05767_ ), .A4(_05770_ ), .ZN(_05771_ ) );
BUF_X4 _20761_ ( .A(_09625_ ), .Z(_05772_ ) );
BUF_X4 _20762_ ( .A(_09121_ ), .Z(_05773_ ) );
AOI22_X1 _20763_ ( .A1(_05772_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_05773_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_05774_ ) );
BUF_X4 _20764_ ( .A(_09552_ ), .Z(_05775_ ) );
BUF_X4 _20765_ ( .A(_09526_ ), .Z(_05776_ ) );
AOI22_X1 _20766_ ( .A1(_05775_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_05776_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05777_ ) );
BUF_X4 _20767_ ( .A(_09081_ ), .Z(_05778_ ) );
NAND3_X1 _20768_ ( .A1(_05774_ ), .A2(_05777_ ), .A3(_05778_ ), .ZN(_05779_ ) );
NAND3_X1 _20769_ ( .A1(_09479_ ), .A2(_05771_ ), .A3(_05779_ ), .ZN(_05780_ ) );
BUF_X4 _20770_ ( .A(_09053_ ), .Z(_05781_ ) );
BUF_X4 _20771_ ( .A(_05740_ ), .Z(_05782_ ) );
BUF_X4 _20772_ ( .A(_09625_ ), .Z(_05783_ ) );
AOI22_X1 _20773_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_05782_ ), .B1(_05783_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05784_ ) );
BUF_X4 _20774_ ( .A(_05737_ ), .Z(_05785_ ) );
AOI22_X1 _20775_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_05773_ ), .B1(_05776_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05786_ ) );
NAND3_X1 _20776_ ( .A1(_05784_ ), .A2(_05785_ ), .A3(_05786_ ), .ZN(_05787_ ) );
AOI22_X1 _20777_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_05782_ ), .B1(_05752_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05788_ ) );
BUF_X4 _20778_ ( .A(_05739_ ), .Z(_05789_ ) );
AOI22_X1 _20779_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_05773_ ), .B1(_05789_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05790_ ) );
NAND3_X1 _20780_ ( .A1(_05788_ ), .A2(_05778_ ), .A3(_05790_ ), .ZN(_05791_ ) );
NAND3_X1 _20781_ ( .A1(_05781_ ), .A2(_05787_ ), .A3(_05791_ ), .ZN(_05792_ ) );
AOI21_X1 _20782_ ( .A(_09115_ ), .B1(_05780_ ), .B2(_05792_ ), .ZN(_05793_ ) );
NOR3_X1 _20783_ ( .A1(_05760_ ), .A2(_08993_ ), .A3(_05793_ ), .ZN(_05794_ ) );
AND3_X1 _20784_ ( .A1(_10428_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_09089_ ), .ZN(_05795_ ) );
AOI221_X4 _20785_ ( .A(_05795_ ), .B1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_05739_ ), .C1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_05740_ ), .ZN(_05796_ ) );
NAND3_X1 _20786_ ( .A1(_09068_ ), .A2(_09092_ ), .A3(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05797_ ) );
NAND3_X1 _20787_ ( .A1(_05796_ ), .A2(_05744_ ), .A3(_05797_ ), .ZN(_05798_ ) );
AND3_X1 _20788_ ( .A1(_10428_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_09089_ ), .ZN(_05799_ ) );
AOI221_X4 _20789_ ( .A(_05799_ ), .B1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_05739_ ), .C1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_05740_ ), .ZN(_05800_ ) );
BUF_X4 _20790_ ( .A(_09081_ ), .Z(_05801_ ) );
NAND3_X1 _20791_ ( .A1(_09068_ ), .A2(_09092_ ), .A3(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05802_ ) );
NAND3_X1 _20792_ ( .A1(_05800_ ), .A2(_05801_ ), .A3(_05802_ ), .ZN(_05803_ ) );
NAND3_X1 _20793_ ( .A1(_05798_ ), .A2(_05803_ ), .A3(_05781_ ), .ZN(_05804_ ) );
OAI211_X1 _20794_ ( .A(_09089_ ), .B(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(_05768_ ), .C2(_05769_ ), .ZN(_05805_ ) );
INV_X1 _20795_ ( .A(_05805_ ), .ZN(_05806_ ) );
AOI221_X4 _20796_ ( .A(_05806_ ), .B1(_05739_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .C2(_09625_ ), .ZN(_05807_ ) );
BUF_X4 _20797_ ( .A(_09067_ ), .Z(_05808_ ) );
BUF_X4 _20798_ ( .A(_05765_ ), .Z(_05809_ ) );
NAND3_X1 _20799_ ( .A1(_05808_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_05809_ ), .ZN(_05810_ ) );
AOI21_X1 _20800_ ( .A(_05751_ ), .B1(_05807_ ), .B2(_05810_ ), .ZN(_05811_ ) );
BUF_X4 _20801_ ( .A(_09121_ ), .Z(_05812_ ) );
AOI22_X1 _20802_ ( .A1(_05782_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_05812_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_05813_ ) );
AOI22_X1 _20803_ ( .A1(_05783_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_05789_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05814_ ) );
AOI21_X1 _20804_ ( .A(_09082_ ), .B1(_05813_ ), .B2(_05814_ ), .ZN(_05815_ ) );
OAI21_X1 _20805_ ( .A(_09479_ ), .B1(_05811_ ), .B2(_05815_ ), .ZN(_05816_ ) );
AOI21_X1 _20806_ ( .A(_09115_ ), .B1(_05804_ ), .B2(_05816_ ), .ZN(_05817_ ) );
AOI22_X1 _20807_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_09552_ ), .B1(_05752_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05818_ ) );
AOI22_X1 _20808_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_05762_ ), .B1(_05789_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05819_ ) );
AOI21_X1 _20809_ ( .A(_09082_ ), .B1(_05818_ ), .B2(_05819_ ), .ZN(_05820_ ) );
AOI22_X1 _20810_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_09552_ ), .B1(_05752_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05821_ ) );
AOI22_X1 _20811_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_05812_ ), .B1(_05789_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05822_ ) );
AOI21_X1 _20812_ ( .A(_05751_ ), .B1(_05821_ ), .B2(_05822_ ), .ZN(_05823_ ) );
OAI21_X1 _20813_ ( .A(_09479_ ), .B1(_05820_ ), .B2(_05823_ ), .ZN(_05824_ ) );
AOI22_X1 _20814_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_05782_ ), .B1(_05752_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05825_ ) );
AOI22_X1 _20815_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_05762_ ), .B1(_05789_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05826_ ) );
NAND3_X1 _20816_ ( .A1(_05825_ ), .A2(_05751_ ), .A3(_05826_ ), .ZN(_05827_ ) );
AOI22_X1 _20817_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_09552_ ), .B1(_05752_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05828_ ) );
AOI22_X1 _20818_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_05762_ ), .B1(_05789_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05829_ ) );
NAND3_X1 _20819_ ( .A1(_05828_ ), .A2(_05778_ ), .A3(_05829_ ), .ZN(_05830_ ) );
NAND3_X1 _20820_ ( .A1(_09053_ ), .A2(_05827_ ), .A3(_05830_ ), .ZN(_05831_ ) );
AOI21_X1 _20821_ ( .A(_09044_ ), .B1(_05824_ ), .B2(_05831_ ), .ZN(_05832_ ) );
NOR3_X1 _20822_ ( .A1(_05817_ ), .A2(_05832_ ), .A3(_08994_ ), .ZN(_05833_ ) );
OAI21_X1 _20823_ ( .A(_09018_ ), .B1(_05794_ ), .B2(_05833_ ), .ZN(_05834_ ) );
AND3_X1 _20824_ ( .A1(_10428_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_05745_ ), .ZN(_05835_ ) );
AOI221_X4 _20825_ ( .A(_05835_ ), .B1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_05739_ ), .C1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_05740_ ), .ZN(_05836_ ) );
NAND3_X1 _20826_ ( .A1(_09068_ ), .A2(_09092_ ), .A3(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05837_ ) );
NAND3_X1 _20827_ ( .A1(_05836_ ), .A2(_09083_ ), .A3(_05837_ ), .ZN(_05838_ ) );
MUX2_X1 _20828_ ( .A(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .S(_05745_ ), .Z(_05839_ ) );
MUX2_X1 _20829_ ( .A(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .S(_05765_ ), .Z(_05840_ ) );
MUX2_X1 _20830_ ( .A(_05839_ ), .B(_05840_ ), .S(_10429_ ), .Z(_05841_ ) );
OAI211_X1 _20831_ ( .A(_05838_ ), .B(_09054_ ), .C1(_09083_ ), .C2(_05841_ ), .ZN(_05842_ ) );
NAND3_X1 _20832_ ( .A1(_09066_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_05745_ ), .ZN(_05843_ ) );
INV_X1 _20833_ ( .A(_05843_ ), .ZN(_05844_ ) );
AOI221_X4 _20834_ ( .A(_05844_ ), .B1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_09121_ ), .C1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_09526_ ), .ZN(_05845_ ) );
NAND3_X1 _20835_ ( .A1(_09068_ ), .A2(_09092_ ), .A3(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05846_ ) );
AOI21_X1 _20836_ ( .A(_05744_ ), .B1(_05845_ ), .B2(_05846_ ), .ZN(_05847_ ) );
BUF_X4 _20837_ ( .A(_09121_ ), .Z(_05848_ ) );
AOI22_X1 _20838_ ( .A1(_05772_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_05848_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_05849_ ) );
AOI22_X1 _20839_ ( .A1(_09553_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_09527_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05850_ ) );
AOI21_X1 _20840_ ( .A(_05801_ ), .B1(_05849_ ), .B2(_05850_ ), .ZN(_05851_ ) );
OAI21_X1 _20841_ ( .A(_09480_ ), .B1(_05847_ ), .B2(_05851_ ), .ZN(_05852_ ) );
NAND3_X1 _20842_ ( .A1(_05842_ ), .A2(_09664_ ), .A3(_05852_ ), .ZN(_05853_ ) );
NAND3_X1 _20843_ ( .A1(_09066_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_05745_ ), .ZN(_05854_ ) );
INV_X1 _20844_ ( .A(_05854_ ), .ZN(_05855_ ) );
AOI221_X4 _20845_ ( .A(_05855_ ), .B1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B2(_09121_ ), .C1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_09526_ ), .ZN(_05856_ ) );
NAND3_X1 _20846_ ( .A1(_09068_ ), .A2(_09092_ ), .A3(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05857_ ) );
AOI21_X1 _20847_ ( .A(_05801_ ), .B1(_05856_ ), .B2(_05857_ ), .ZN(_05858_ ) );
NAND3_X1 _20848_ ( .A1(_09066_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_05745_ ), .ZN(_05859_ ) );
INV_X1 _20849_ ( .A(_05859_ ), .ZN(_05860_ ) );
AOI221_X4 _20850_ ( .A(_05860_ ), .B1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_09121_ ), .C1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_09526_ ), .ZN(_05861_ ) );
NAND3_X1 _20851_ ( .A1(_09068_ ), .A2(_09092_ ), .A3(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05862_ ) );
AOI21_X1 _20852_ ( .A(_05785_ ), .B1(_05861_ ), .B2(_05862_ ), .ZN(_05863_ ) );
OAI21_X1 _20853_ ( .A(_09480_ ), .B1(_05858_ ), .B2(_05863_ ), .ZN(_05864_ ) );
BUF_X4 _20854_ ( .A(_09526_ ), .Z(_05865_ ) );
AOI22_X1 _20855_ ( .A1(_05772_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_05865_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05866_ ) );
NAND3_X1 _20856_ ( .A1(_09068_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_05809_ ), .ZN(_05867_ ) );
BUF_X4 _20857_ ( .A(_05768_ ), .Z(_05868_ ) );
BUF_X4 _20858_ ( .A(_05769_ ), .Z(_05869_ ) );
OAI211_X1 _20859_ ( .A(_05766_ ), .B(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C1(_05868_ ), .C2(_05869_ ), .ZN(_05870_ ) );
NAND4_X1 _20860_ ( .A1(_05866_ ), .A2(_05744_ ), .A3(_05867_ ), .A4(_05870_ ), .ZN(_05871_ ) );
AOI22_X1 _20861_ ( .A1(_09553_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_05848_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_05872_ ) );
AOI22_X1 _20862_ ( .A1(_09626_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_05865_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05873_ ) );
NAND3_X1 _20863_ ( .A1(_05872_ ), .A2(_05873_ ), .A3(_05801_ ), .ZN(_05874_ ) );
NAND3_X1 _20864_ ( .A1(_09054_ ), .A2(_05871_ ), .A3(_05874_ ), .ZN(_05875_ ) );
NAND3_X1 _20865_ ( .A1(_05864_ ), .A2(_09045_ ), .A3(_05875_ ), .ZN(_05876_ ) );
NAND3_X1 _20866_ ( .A1(_05853_ ), .A2(_08995_ ), .A3(_05876_ ), .ZN(_05877_ ) );
NAND3_X1 _20867_ ( .A1(_09066_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_09089_ ), .ZN(_05878_ ) );
INV_X1 _20868_ ( .A(_05878_ ), .ZN(_05879_ ) );
AOI221_X4 _20869_ ( .A(_05879_ ), .B1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_09120_ ), .C1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_09526_ ), .ZN(_05880_ ) );
NAND3_X1 _20870_ ( .A1(_05808_ ), .A2(_09092_ ), .A3(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05881_ ) );
AOI21_X1 _20871_ ( .A(_05785_ ), .B1(_05880_ ), .B2(_05881_ ), .ZN(_05882_ ) );
AOI22_X1 _20872_ ( .A1(_05775_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_05762_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_05883_ ) );
AOI22_X1 _20873_ ( .A1(_05761_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_05776_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05884_ ) );
AOI21_X1 _20874_ ( .A(_09082_ ), .B1(_05883_ ), .B2(_05884_ ), .ZN(_05885_ ) );
OAI21_X1 _20875_ ( .A(_09480_ ), .B1(_05882_ ), .B2(_05885_ ), .ZN(_05886_ ) );
AND3_X1 _20876_ ( .A1(_05748_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_05765_ ), .ZN(_05887_ ) );
OAI211_X1 _20877_ ( .A(_09090_ ), .B(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_05768_ ), .C2(_05769_ ), .ZN(_05888_ ) );
NAND3_X1 _20878_ ( .A1(_09067_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_05765_ ), .ZN(_05889_ ) );
NAND2_X1 _20879_ ( .A1(_05888_ ), .A2(_05889_ ), .ZN(_05890_ ) );
AND3_X1 _20880_ ( .A1(_09067_ ), .A2(_09090_ ), .A3(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05891_ ) );
NOR3_X1 _20881_ ( .A1(_05887_ ), .A2(_05890_ ), .A3(_05891_ ), .ZN(_05892_ ) );
AOI22_X1 _20882_ ( .A1(_05740_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_09526_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05893_ ) );
NAND3_X1 _20883_ ( .A1(_05748_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_05765_ ), .ZN(_05894_ ) );
NAND3_X1 _20884_ ( .A1(_09067_ ), .A2(_09091_ ), .A3(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05895_ ) );
AND3_X1 _20885_ ( .A1(_05893_ ), .A2(_05894_ ), .A3(_05895_ ), .ZN(_05896_ ) );
MUX2_X1 _20886_ ( .A(_05892_ ), .B(_05896_ ), .S(_09082_ ), .Z(_05897_ ) );
OAI211_X1 _20887_ ( .A(_05886_ ), .B(_09045_ ), .C1(_09480_ ), .C2(_05897_ ), .ZN(_05898_ ) );
AOI22_X1 _20888_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_09553_ ), .B1(_05772_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05899_ ) );
AOI22_X1 _20889_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_05848_ ), .B1(_05865_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05900_ ) );
NAND3_X1 _20890_ ( .A1(_05899_ ), .A2(_09083_ ), .A3(_05900_ ), .ZN(_05901_ ) );
AOI22_X1 _20891_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_09553_ ), .B1(_05772_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05902_ ) );
AOI22_X1 _20892_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_05848_ ), .B1(_05865_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05903_ ) );
NAND3_X1 _20893_ ( .A1(_05902_ ), .A2(_05744_ ), .A3(_05903_ ), .ZN(_05904_ ) );
NAND3_X1 _20894_ ( .A1(_09480_ ), .A2(_05901_ ), .A3(_05904_ ), .ZN(_05905_ ) );
AOI22_X1 _20895_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_09553_ ), .B1(_05772_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05906_ ) );
AOI22_X1 _20896_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_05848_ ), .B1(_09527_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05907_ ) );
NAND3_X1 _20897_ ( .A1(_05906_ ), .A2(_05744_ ), .A3(_05907_ ), .ZN(_05908_ ) );
AOI22_X1 _20898_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_09553_ ), .B1(_05772_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05909_ ) );
AOI22_X1 _20899_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_05848_ ), .B1(_09527_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05910_ ) );
NAND3_X1 _20900_ ( .A1(_05909_ ), .A2(_05801_ ), .A3(_05910_ ), .ZN(_05911_ ) );
NAND3_X1 _20901_ ( .A1(_09054_ ), .A2(_05908_ ), .A3(_05911_ ), .ZN(_05912_ ) );
NAND3_X1 _20902_ ( .A1(_05905_ ), .A2(_09664_ ), .A3(_05912_ ), .ZN(_05913_ ) );
NAND3_X1 _20903_ ( .A1(_05898_ ), .A2(_08993_ ), .A3(_05913_ ), .ZN(_05914_ ) );
NAND3_X1 _20904_ ( .A1(_05877_ ), .A2(_05914_ ), .A3(_09019_ ), .ZN(_05915_ ) );
AND3_X1 _20905_ ( .A1(_05834_ ), .A2(_09034_ ), .A3(_05915_ ), .ZN(_05916_ ) );
AND3_X1 _20906_ ( .A1(_10428_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_09089_ ), .ZN(_05917_ ) );
AOI221_X1 _20907_ ( .A(_05917_ ), .B1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_05739_ ), .C1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_05740_ ), .ZN(_05918_ ) );
NAND3_X1 _20908_ ( .A1(_05808_ ), .A2(_09092_ ), .A3(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05919_ ) );
NAND3_X1 _20909_ ( .A1(_05918_ ), .A2(_05778_ ), .A3(_05919_ ), .ZN(_05920_ ) );
MUX2_X1 _20910_ ( .A(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .S(_05745_ ), .Z(_05921_ ) );
MUX2_X1 _20911_ ( .A(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .S(_05745_ ), .Z(_05922_ ) );
MUX2_X1 _20912_ ( .A(_05921_ ), .B(_05922_ ), .S(_05748_ ), .Z(_05923_ ) );
OAI211_X1 _20913_ ( .A(_05920_ ), .B(_09479_ ), .C1(_09083_ ), .C2(_05923_ ), .ZN(_05924_ ) );
AOI22_X1 _20914_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_05775_ ), .B1(_05783_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05925_ ) );
AOI22_X1 _20915_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_05773_ ), .B1(_05776_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05926_ ) );
NAND3_X1 _20916_ ( .A1(_05925_ ), .A2(_05801_ ), .A3(_05926_ ), .ZN(_05927_ ) );
AOI22_X1 _20917_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_05775_ ), .B1(_05783_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05928_ ) );
AOI22_X1 _20918_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_05773_ ), .B1(_05776_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05929_ ) );
NAND3_X1 _20919_ ( .A1(_05928_ ), .A2(_05785_ ), .A3(_05929_ ), .ZN(_05930_ ) );
NAND3_X1 _20920_ ( .A1(_05781_ ), .A2(_05927_ ), .A3(_05930_ ), .ZN(_05931_ ) );
AOI21_X1 _20921_ ( .A(_09045_ ), .B1(_05924_ ), .B2(_05931_ ), .ZN(_05932_ ) );
AOI22_X1 _20922_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_05775_ ), .B1(_05783_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05933_ ) );
AOI22_X1 _20923_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_05773_ ), .B1(_05776_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05934_ ) );
NAND3_X1 _20924_ ( .A1(_05933_ ), .A2(_05785_ ), .A3(_05934_ ), .ZN(_05935_ ) );
AOI22_X1 _20925_ ( .A1(_05782_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_05812_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_05936_ ) );
BUF_X4 _20926_ ( .A(_09090_ ), .Z(_05937_ ) );
NAND3_X1 _20927_ ( .A1(_05764_ ), .A2(_05937_ ), .A3(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05938_ ) );
OAI211_X1 _20928_ ( .A(_09091_ ), .B(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_05768_ ), .C2(_05769_ ), .ZN(_05939_ ) );
NAND4_X1 _20929_ ( .A1(_05936_ ), .A2(_05778_ ), .A3(_05938_ ), .A4(_05939_ ), .ZN(_05940_ ) );
NAND3_X1 _20930_ ( .A1(_09479_ ), .A2(_05935_ ), .A3(_05940_ ), .ZN(_05941_ ) );
AOI22_X1 _20931_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_05782_ ), .B1(_05752_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05942_ ) );
AOI22_X1 _20932_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_05773_ ), .B1(_05789_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05943_ ) );
NAND3_X1 _20933_ ( .A1(_05942_ ), .A2(_05785_ ), .A3(_05943_ ), .ZN(_05944_ ) );
AOI22_X1 _20934_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_09552_ ), .B1(_05752_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05945_ ) );
AOI22_X1 _20935_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_05762_ ), .B1(_05789_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05946_ ) );
NAND3_X1 _20936_ ( .A1(_05945_ ), .A2(_05778_ ), .A3(_05946_ ), .ZN(_05947_ ) );
NAND3_X1 _20937_ ( .A1(_05781_ ), .A2(_05944_ ), .A3(_05947_ ), .ZN(_05948_ ) );
AOI21_X1 _20938_ ( .A(_09115_ ), .B1(_05941_ ), .B2(_05948_ ), .ZN(_05949_ ) );
OAI21_X1 _20939_ ( .A(_08994_ ), .B1(_05932_ ), .B2(_05949_ ), .ZN(_05950_ ) );
AOI22_X1 _20940_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_05782_ ), .B1(_05783_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05951_ ) );
AOI22_X1 _20941_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_05773_ ), .B1(_05776_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05952_ ) );
NAND3_X1 _20942_ ( .A1(_05951_ ), .A2(_05778_ ), .A3(_05952_ ), .ZN(_05953_ ) );
AOI22_X1 _20943_ ( .A1(_05775_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_05762_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_05954_ ) );
AOI22_X1 _20944_ ( .A1(_05761_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_05776_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05955_ ) );
NAND3_X1 _20945_ ( .A1(_05954_ ), .A2(_05955_ ), .A3(_05785_ ), .ZN(_05956_ ) );
NAND3_X1 _20946_ ( .A1(_05781_ ), .A2(_05953_ ), .A3(_05956_ ), .ZN(_05957_ ) );
AOI22_X1 _20947_ ( .A1(_05740_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_05739_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05958_ ) );
NAND3_X1 _20948_ ( .A1(_09067_ ), .A2(_09090_ ), .A3(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05959_ ) );
NAND3_X1 _20949_ ( .A1(_05748_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_05765_ ), .ZN(_05960_ ) );
AND3_X1 _20950_ ( .A1(_05958_ ), .A2(_05959_ ), .A3(_05960_ ), .ZN(_05961_ ) );
AOI22_X1 _20951_ ( .A1(_05740_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_05739_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05962_ ) );
NAND3_X1 _20952_ ( .A1(_09067_ ), .A2(_09090_ ), .A3(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05963_ ) );
NAND3_X1 _20953_ ( .A1(_05748_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_05765_ ), .ZN(_05964_ ) );
AND3_X1 _20954_ ( .A1(_05962_ ), .A2(_05963_ ), .A3(_05964_ ), .ZN(_05965_ ) );
MUX2_X1 _20955_ ( .A(_05961_ ), .B(_05965_ ), .S(_09082_ ), .Z(_05966_ ) );
OAI211_X1 _20956_ ( .A(_09045_ ), .B(_05957_ ), .C1(_05966_ ), .C2(_09054_ ), .ZN(_05967_ ) );
AOI22_X1 _20957_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_09553_ ), .B1(_05761_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05968_ ) );
AOI22_X1 _20958_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_05848_ ), .B1(_09527_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05969_ ) );
NAND3_X1 _20959_ ( .A1(_05968_ ), .A2(_05744_ ), .A3(_05969_ ), .ZN(_05970_ ) );
AOI22_X1 _20960_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_05775_ ), .B1(_05761_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05971_ ) );
AOI22_X1 _20961_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_05848_ ), .B1(_09527_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05972_ ) );
NAND3_X1 _20962_ ( .A1(_05971_ ), .A2(_05801_ ), .A3(_05972_ ), .ZN(_05973_ ) );
NAND3_X1 _20963_ ( .A1(_09480_ ), .A2(_05970_ ), .A3(_05973_ ), .ZN(_05974_ ) );
AOI22_X1 _20964_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_05782_ ), .B1(_05783_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05975_ ) );
AOI22_X1 _20965_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_05773_ ), .B1(_05776_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05976_ ) );
AOI21_X1 _20966_ ( .A(_09082_ ), .B1(_05975_ ), .B2(_05976_ ), .ZN(_05977_ ) );
AOI22_X1 _20967_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_09552_ ), .B1(_05752_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05978_ ) );
AOI22_X1 _20968_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_05812_ ), .B1(_05789_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05979_ ) );
AOI21_X1 _20969_ ( .A(_05751_ ), .B1(_05978_ ), .B2(_05979_ ), .ZN(_05980_ ) );
OAI21_X1 _20970_ ( .A(_05781_ ), .B1(_05977_ ), .B2(_05980_ ), .ZN(_05981_ ) );
NAND3_X1 _20971_ ( .A1(_05974_ ), .A2(_09664_ ), .A3(_05981_ ), .ZN(_05982_ ) );
NAND3_X1 _20972_ ( .A1(_05967_ ), .A2(_05982_ ), .A3(_08993_ ), .ZN(_05983_ ) );
AOI21_X1 _20973_ ( .A(_09019_ ), .B1(_05950_ ), .B2(_05983_ ), .ZN(_05984_ ) );
AND3_X1 _20974_ ( .A1(_10428_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_09089_ ), .ZN(_05985_ ) );
AOI221_X1 _20975_ ( .A(_05985_ ), .B1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_05739_ ), .C1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_05740_ ), .ZN(_05986_ ) );
NAND3_X1 _20976_ ( .A1(_05808_ ), .A2(_09092_ ), .A3(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05987_ ) );
NAND3_X1 _20977_ ( .A1(_05986_ ), .A2(_05801_ ), .A3(_05987_ ), .ZN(_05988_ ) );
AOI22_X1 _20978_ ( .A1(_05775_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_05776_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05989_ ) );
OAI211_X1 _20979_ ( .A(_05766_ ), .B(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C1(_05868_ ), .C2(_05869_ ), .ZN(_05990_ ) );
NAND3_X1 _20980_ ( .A1(_05808_ ), .A2(_05937_ ), .A3(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05991_ ) );
NAND3_X1 _20981_ ( .A1(_05989_ ), .A2(_05990_ ), .A3(_05991_ ), .ZN(_05992_ ) );
OAI211_X1 _20982_ ( .A(_05988_ ), .B(_09479_ ), .C1(_09083_ ), .C2(_05992_ ), .ZN(_05993_ ) );
AOI22_X1 _20983_ ( .A1(_05775_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_09527_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05994_ ) );
OAI211_X1 _20984_ ( .A(_05766_ ), .B(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C1(_05868_ ), .C2(_05869_ ), .ZN(_05995_ ) );
NAND3_X1 _20985_ ( .A1(_05808_ ), .A2(_05937_ ), .A3(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05996_ ) );
NAND4_X1 _20986_ ( .A1(_05994_ ), .A2(_05785_ ), .A3(_05995_ ), .A4(_05996_ ), .ZN(_05997_ ) );
AOI22_X1 _20987_ ( .A1(_09553_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_05773_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_05998_ ) );
AOI22_X1 _20988_ ( .A1(_05772_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_09527_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05999_ ) );
NAND3_X1 _20989_ ( .A1(_05998_ ), .A2(_05999_ ), .A3(_05801_ ), .ZN(_06000_ ) );
NAND3_X1 _20990_ ( .A1(_05781_ ), .A2(_05997_ ), .A3(_06000_ ), .ZN(_06001_ ) );
NAND3_X1 _20991_ ( .A1(_05993_ ), .A2(_09045_ ), .A3(_06001_ ), .ZN(_06002_ ) );
AOI22_X1 _20992_ ( .A1(_05772_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_05762_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06003_ ) );
OAI211_X1 _20993_ ( .A(_05937_ ), .B(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_05868_ ), .C2(_05869_ ), .ZN(_06004_ ) );
NAND3_X1 _20994_ ( .A1(_05808_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_05766_ ), .ZN(_06005_ ) );
NAND4_X1 _20995_ ( .A1(_06003_ ), .A2(_05785_ ), .A3(_06004_ ), .A4(_06005_ ), .ZN(_06006_ ) );
AOI22_X1 _20996_ ( .A1(_05772_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_05762_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06007_ ) );
OAI211_X1 _20997_ ( .A(_05937_ ), .B(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_05868_ ), .C2(_05869_ ), .ZN(_06008_ ) );
NAND3_X1 _20998_ ( .A1(_05808_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_05766_ ), .ZN(_06009_ ) );
NAND4_X1 _20999_ ( .A1(_06007_ ), .A2(_05778_ ), .A3(_06008_ ), .A4(_06009_ ), .ZN(_06010_ ) );
NAND3_X1 _21000_ ( .A1(_09480_ ), .A2(_06006_ ), .A3(_06010_ ), .ZN(_06011_ ) );
AOI22_X1 _21001_ ( .A1(_05761_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_05812_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06012_ ) );
OAI211_X1 _21002_ ( .A(_09091_ ), .B(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_05768_ ), .C2(_05769_ ), .ZN(_06013_ ) );
NAND3_X1 _21003_ ( .A1(_05764_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_05766_ ), .ZN(_06014_ ) );
NAND4_X1 _21004_ ( .A1(_06012_ ), .A2(_05751_ ), .A3(_06013_ ), .A4(_06014_ ), .ZN(_06015_ ) );
AOI22_X1 _21005_ ( .A1(_05783_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_05812_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06016_ ) );
OAI211_X1 _21006_ ( .A(_09091_ ), .B(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_05768_ ), .C2(_05769_ ), .ZN(_06017_ ) );
BUF_X4 _21007_ ( .A(_05765_ ), .Z(_06018_ ) );
NAND3_X1 _21008_ ( .A1(_05764_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06018_ ), .ZN(_06019_ ) );
NAND4_X1 _21009_ ( .A1(_06016_ ), .A2(_09082_ ), .A3(_06017_ ), .A4(_06019_ ), .ZN(_06020_ ) );
NAND3_X1 _21010_ ( .A1(_05781_ ), .A2(_06015_ ), .A3(_06020_ ), .ZN(_06021_ ) );
NAND3_X1 _21011_ ( .A1(_06011_ ), .A2(_09115_ ), .A3(_06021_ ), .ZN(_06022_ ) );
NAND3_X1 _21012_ ( .A1(_06002_ ), .A2(_08994_ ), .A3(_06022_ ), .ZN(_06023_ ) );
AOI22_X1 _21013_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_05775_ ), .B1(_05761_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06024_ ) );
AOI22_X1 _21014_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_05848_ ), .B1(_09527_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06025_ ) );
NAND3_X1 _21015_ ( .A1(_06024_ ), .A2(_05785_ ), .A3(_06025_ ), .ZN(_06026_ ) );
AOI22_X1 _21016_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_05848_ ), .B1(_09527_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06027_ ) );
AOI22_X1 _21017_ ( .A1(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_05782_ ), .B1(_05783_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06028_ ) );
NAND3_X1 _21018_ ( .A1(_06027_ ), .A2(_05801_ ), .A3(_06028_ ), .ZN(_06029_ ) );
NAND3_X1 _21019_ ( .A1(_09480_ ), .A2(_06026_ ), .A3(_06029_ ), .ZN(_06030_ ) );
AOI22_X1 _21020_ ( .A1(_05761_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_05812_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06031_ ) );
OAI211_X1 _21021_ ( .A(_05937_ ), .B(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_05868_ ), .C2(_05869_ ), .ZN(_06032_ ) );
NAND3_X1 _21022_ ( .A1(_05764_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_05766_ ), .ZN(_06033_ ) );
NAND4_X1 _21023_ ( .A1(_06031_ ), .A2(_05778_ ), .A3(_06032_ ), .A4(_06033_ ), .ZN(_06034_ ) );
AOI22_X1 _21024_ ( .A1(_05761_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_05812_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06035_ ) );
OAI211_X1 _21025_ ( .A(_09091_ ), .B(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_05768_ ), .C2(_05769_ ), .ZN(_06036_ ) );
NAND3_X1 _21026_ ( .A1(_05764_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06018_ ), .ZN(_06037_ ) );
NAND4_X1 _21027_ ( .A1(_06035_ ), .A2(_05751_ ), .A3(_06036_ ), .A4(_06037_ ), .ZN(_06038_ ) );
NAND3_X1 _21028_ ( .A1(_05781_ ), .A2(_06034_ ), .A3(_06038_ ), .ZN(_06039_ ) );
NAND3_X1 _21029_ ( .A1(_06030_ ), .A2(_09664_ ), .A3(_06039_ ), .ZN(_06040_ ) );
AOI22_X1 _21030_ ( .A1(_05761_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_05762_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06041_ ) );
NAND3_X1 _21031_ ( .A1(_05808_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_05766_ ), .ZN(_06042_ ) );
OAI211_X1 _21032_ ( .A(_05937_ ), .B(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_05768_ ), .C2(_05769_ ), .ZN(_06043_ ) );
NAND4_X1 _21033_ ( .A1(_06041_ ), .A2(_05751_ ), .A3(_06042_ ), .A4(_06043_ ), .ZN(_06044_ ) );
AOI22_X1 _21034_ ( .A1(_05782_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_05812_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06045_ ) );
NAND3_X1 _21035_ ( .A1(_05764_ ), .A2(_05937_ ), .A3(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06046_ ) );
OAI211_X1 _21036_ ( .A(_09091_ ), .B(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_05768_ ), .C2(_05769_ ), .ZN(_06047_ ) );
NAND4_X1 _21037_ ( .A1(_06045_ ), .A2(_05778_ ), .A3(_06046_ ), .A4(_06047_ ), .ZN(_06048_ ) );
NAND3_X1 _21038_ ( .A1(_09480_ ), .A2(_06044_ ), .A3(_06048_ ), .ZN(_06049_ ) );
AOI22_X1 _21039_ ( .A1(_05783_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_05812_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06050_ ) );
NAND3_X1 _21040_ ( .A1(_05764_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06018_ ), .ZN(_06051_ ) );
NAND3_X1 _21041_ ( .A1(_10429_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_05937_ ), .ZN(_06052_ ) );
NAND4_X1 _21042_ ( .A1(_06050_ ), .A2(_05751_ ), .A3(_06051_ ), .A4(_06052_ ), .ZN(_06053_ ) );
AOI22_X1 _21043_ ( .A1(_09552_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_05789_ ), .B2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06054_ ) );
NAND3_X1 _21044_ ( .A1(_05764_ ), .A2(_05937_ ), .A3(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06055_ ) );
NAND3_X1 _21045_ ( .A1(_10429_ ), .A2(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06018_ ), .ZN(_06056_ ) );
NAND4_X1 _21046_ ( .A1(_06054_ ), .A2(_09082_ ), .A3(_06055_ ), .A4(_06056_ ), .ZN(_06057_ ) );
NAND3_X1 _21047_ ( .A1(_05781_ ), .A2(_06053_ ), .A3(_06057_ ), .ZN(_06058_ ) );
NAND3_X1 _21048_ ( .A1(_06049_ ), .A2(_09045_ ), .A3(_06058_ ), .ZN(_06059_ ) );
NAND3_X1 _21049_ ( .A1(_06040_ ), .A2(_06059_ ), .A3(_08993_ ), .ZN(_06060_ ) );
AOI21_X1 _21050_ ( .A(_09018_ ), .B1(_06023_ ), .B2(_06060_ ), .ZN(_06061_ ) );
OAI21_X1 _21051_ ( .A(_09138_ ), .B1(_05984_ ), .B2(_06061_ ), .ZN(_06062_ ) );
NAND2_X1 _21052_ ( .A1(_06062_ ), .A2(_05734_ ), .ZN(_06063_ ) );
NOR2_X4 _21053_ ( .A1(_05916_ ), .A2(_06063_ ), .ZN(\load_data_out[10] ) );
NOR2_X4 _21054_ ( .A1(\load_data_out[10] ), .A2(_05735_ ), .ZN(_06064_ ) );
NOR2_X2 _21055_ ( .A1(_06064_ ), .A2(_08944_ ), .ZN(_06065_ ) );
AOI21_X1 _21056_ ( .A(_05732_ ), .B1(_05736_ ), .B2(_06065_ ), .ZN(_06066_ ) );
AOI21_X1 _21057_ ( .A(_08914_ ), .B1(_08921_ ), .B2(\ifu_rdata[2] ), .ZN(_06067_ ) );
AOI21_X1 _21058_ ( .A(fanout_net_75 ), .B1(_05730_ ), .B2(_06067_ ), .ZN(_06068_ ) );
INV_X1 _21059_ ( .A(\ifu_rdata[7] ), .ZN(_06069_ ) );
INV_X1 _21060_ ( .A(\ifu_rdata[8] ), .ZN(_06070_ ) );
NAND3_X1 _21061_ ( .A1(_06069_ ), .A2(_06070_ ), .A3(alu_result_out_$_XNOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B_$_OR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_06071_ ) );
AND3_X1 _21062_ ( .A1(_06068_ ), .A2(_08586_ ), .A3(_06071_ ), .ZN(_06072_ ) );
NOR2_X1 _21063_ ( .A1(_06069_ ), .A2(\ifu_rdata[8] ), .ZN(_06073_ ) );
NAND2_X2 _21064_ ( .A1(_06072_ ), .A2(_06073_ ), .ZN(_06074_ ) );
BUF_X4 _21065_ ( .A(_06074_ ), .Z(_06075_ ) );
NOR2_X1 _21066_ ( .A1(_06066_ ), .A2(_06075_ ), .ZN(_00005_ ) );
BUF_X4 _21067_ ( .A(_06074_ ), .Z(_06076_ ) );
BUF_X2 _21068_ ( .A(_05734_ ), .Z(_06077_ ) );
INV_X1 _21069_ ( .A(_08913_ ), .ZN(_06078_ ) );
AND2_X1 _21070_ ( .A1(\alu_result_out[30] ), .A2(_06078_ ), .ZN(_06079_ ) );
OAI21_X1 _21071_ ( .A(_06065_ ), .B1(_06077_ ), .B2(_06079_ ), .ZN(_06080_ ) );
BUF_X4 _21072_ ( .A(_05729_ ), .Z(_06081_ ) );
BUF_X4 _21073_ ( .A(_08908_ ), .Z(_06082_ ) );
AOI22_X1 _21074_ ( .A1(\alu_result_out[30] ), .A2(_06081_ ), .B1(_06082_ ), .B2(_09305_ ), .ZN(_06083_ ) );
AOI21_X1 _21075_ ( .A(_06076_ ), .B1(_06080_ ), .B2(_06083_ ), .ZN(_00006_ ) );
NOR2_X1 _21076_ ( .A1(_09425_ ), .A2(_09105_ ), .ZN(_06084_ ) );
NOR3_X1 _21077_ ( .A1(_08910_ ), .A2(\ifu_rdata[2] ), .A3(\ifu_rdata[5] ), .ZN(_06085_ ) );
AND2_X1 _21078_ ( .A1(_06085_ ), .A2(_08902_ ), .ZN(_06086_ ) );
OR2_X1 _21079_ ( .A1(_05729_ ), .A2(_06086_ ), .ZN(_06087_ ) );
BUF_X2 _21080_ ( .A(_06087_ ), .Z(_06088_ ) );
AND2_X1 _21081_ ( .A1(\alu_result_out[21] ), .A2(_06088_ ), .ZN(_06089_ ) );
NOR3_X1 _21082_ ( .A1(\load_data_out[10] ), .A2(_06084_ ), .A3(_06089_ ), .ZN(_06090_ ) );
NOR2_X1 _21083_ ( .A1(_06090_ ), .A2(_06075_ ), .ZN(_00007_ ) );
INV_X1 _21084_ ( .A(\load_data_out[10] ), .ZN(_06091_ ) );
BUF_X4 _21085_ ( .A(_06091_ ), .Z(_06092_ ) );
AOI22_X1 _21086_ ( .A1(\alu_result_out[20] ), .A2(_06088_ ), .B1(_06082_ ), .B2(_09320_ ), .ZN(_06093_ ) );
AOI21_X1 _21087_ ( .A(_06076_ ), .B1(_06092_ ), .B2(_06093_ ), .ZN(_00008_ ) );
NOR2_X1 _21088_ ( .A1(_09329_ ), .A2(_09105_ ), .ZN(_06094_ ) );
AND2_X1 _21089_ ( .A1(\alu_result_out[19] ), .A2(_06088_ ), .ZN(_06095_ ) );
NOR3_X1 _21090_ ( .A1(\load_data_out[10] ), .A2(_06094_ ), .A3(_06095_ ), .ZN(_06096_ ) );
NOR2_X1 _21091_ ( .A1(_06096_ ), .A2(_06075_ ), .ZN(_00009_ ) );
AOI22_X1 _21092_ ( .A1(\alu_result_out[18] ), .A2(_06088_ ), .B1(_06082_ ), .B2(_09331_ ), .ZN(_06097_ ) );
AOI21_X1 _21093_ ( .A(_06076_ ), .B1(_06092_ ), .B2(_06097_ ), .ZN(_00010_ ) );
NOR2_X1 _21094_ ( .A1(_09340_ ), .A2(_09105_ ), .ZN(_06098_ ) );
AND2_X1 _21095_ ( .A1(\alu_result_out[17] ), .A2(_06087_ ), .ZN(_06099_ ) );
NOR3_X1 _21096_ ( .A1(\load_data_out[10] ), .A2(_06098_ ), .A3(_06099_ ), .ZN(_06100_ ) );
NOR2_X1 _21097_ ( .A1(_06100_ ), .A2(_06075_ ), .ZN(_00011_ ) );
INV_X1 _21098_ ( .A(_08944_ ), .ZN(_06101_ ) );
BUF_X4 _21099_ ( .A(_06101_ ), .Z(_06102_ ) );
AND3_X1 _21100_ ( .A1(\alu_result_out[16] ), .A2(_06078_ ), .A3(_05735_ ), .ZN(_06103_ ) );
OAI21_X1 _21101_ ( .A(_06102_ ), .B1(\load_data_out[10] ), .B2(_06103_ ), .ZN(_06104_ ) );
AOI22_X1 _21102_ ( .A1(\alu_result_out[16] ), .A2(_06081_ ), .B1(_06082_ ), .B2(_09343_ ), .ZN(_06105_ ) );
AOI21_X1 _21103_ ( .A(_06076_ ), .B1(_06104_ ), .B2(_06105_ ), .ZN(_00012_ ) );
AND2_X1 _21104_ ( .A1(\alu_result_out[15] ), .A2(_06078_ ), .ZN(_06106_ ) );
OAI21_X1 _21105_ ( .A(_06065_ ), .B1(_06077_ ), .B2(_06106_ ), .ZN(_06107_ ) );
NAND2_X1 _21106_ ( .A1(\alu_result_out[15] ), .A2(_06081_ ), .ZN(_06108_ ) );
OR2_X1 _21107_ ( .A1(_09354_ ), .A2(_08928_ ), .ZN(_06109_ ) );
AND3_X2 _21108_ ( .A1(_06107_ ), .A2(_06108_ ), .A3(_06109_ ), .ZN(_06110_ ) );
NOR2_X1 _21109_ ( .A1(_06110_ ), .A2(_06075_ ), .ZN(_00013_ ) );
AOI22_X1 _21110_ ( .A1(\alu_result_out[14] ), .A2(_06088_ ), .B1(_06082_ ), .B2(_09357_ ), .ZN(_06111_ ) );
AOI21_X1 _21111_ ( .A(_06076_ ), .B1(_06092_ ), .B2(_06111_ ), .ZN(_00014_ ) );
AOI22_X1 _21112_ ( .A1(\alu_result_out[13] ), .A2(_06088_ ), .B1(_06082_ ), .B2(_09364_ ), .ZN(_06112_ ) );
AOI21_X1 _21113_ ( .A(_06076_ ), .B1(_06092_ ), .B2(_06112_ ), .ZN(_00015_ ) );
AND3_X1 _21114_ ( .A1(\alu_result_out[12] ), .A2(_06078_ ), .A3(_05735_ ), .ZN(_06113_ ) );
OAI21_X1 _21115_ ( .A(_06102_ ), .B1(\load_data_out[10] ), .B2(_06113_ ), .ZN(_06114_ ) );
AOI22_X1 _21116_ ( .A1(\alu_result_out[12] ), .A2(_06081_ ), .B1(_06082_ ), .B2(_09368_ ), .ZN(_06115_ ) );
AOI21_X1 _21117_ ( .A(_06076_ ), .B1(_06114_ ), .B2(_06115_ ), .ZN(_00016_ ) );
AND2_X1 _21118_ ( .A1(\alu_result_out[29] ), .A2(_06078_ ), .ZN(_06116_ ) );
OAI21_X1 _21119_ ( .A(_06065_ ), .B1(_06077_ ), .B2(_06116_ ), .ZN(_06117_ ) );
NAND2_X1 _21120_ ( .A1(\alu_result_out[29] ), .A2(_06081_ ), .ZN(_06118_ ) );
OR2_X1 _21121_ ( .A1(_09315_ ), .A2(_08928_ ), .ZN(_06119_ ) );
AND3_X2 _21122_ ( .A1(_06117_ ), .A2(_06118_ ), .A3(_06119_ ), .ZN(_06120_ ) );
NOR2_X1 _21123_ ( .A1(_06120_ ), .A2(_06075_ ), .ZN(_00017_ ) );
NOR2_X1 _21124_ ( .A1(_09376_ ), .A2(_09105_ ), .ZN(_06121_ ) );
AND2_X1 _21125_ ( .A1(\alu_result_out[11] ), .A2(_06087_ ), .ZN(_06122_ ) );
NOR3_X1 _21126_ ( .A1(\load_data_out[10] ), .A2(_06121_ ), .A3(_06122_ ), .ZN(_06123_ ) );
NOR2_X1 _21127_ ( .A1(_06123_ ), .A2(_06075_ ), .ZN(_00018_ ) );
AND3_X1 _21128_ ( .A1(\alu_result_out[10] ), .A2(_06078_ ), .A3(_05735_ ), .ZN(_06124_ ) );
OAI21_X1 _21129_ ( .A(_06101_ ), .B1(\load_data_out[10] ), .B2(_06124_ ), .ZN(_06125_ ) );
NAND2_X1 _21130_ ( .A1(\alu_result_out[10] ), .A2(_06081_ ), .ZN(_06126_ ) );
OR3_X1 _21131_ ( .A1(_08928_ ), .A2(_09375_ ), .A3(_09382_ ), .ZN(_06127_ ) );
AND3_X1 _21132_ ( .A1(_06125_ ), .A2(_06126_ ), .A3(_06127_ ), .ZN(_06128_ ) );
NOR2_X1 _21133_ ( .A1(_06128_ ), .A2(_06075_ ), .ZN(_00019_ ) );
OAI22_X1 _21134_ ( .A1(_10070_ ), .A2(_05731_ ), .B1(_09105_ ), .B2(_09040_ ), .ZN(_06129_ ) );
OR2_X2 _21135_ ( .A1(_08913_ ), .A2(_05734_ ), .ZN(_06130_ ) );
OAI22_X1 _21136_ ( .A1(_05916_ ), .A2(_06063_ ), .B1(_10012_ ), .B2(_06130_ ), .ZN(_06131_ ) );
AOI21_X1 _21137_ ( .A(_06129_ ), .B1(_06131_ ), .B2(_06102_ ), .ZN(_06132_ ) );
NOR2_X1 _21138_ ( .A1(_06132_ ), .A2(_06075_ ), .ZN(_00020_ ) );
NAND2_X1 _21139_ ( .A1(_09023_ ), .A2(_08908_ ), .ZN(_06133_ ) );
OAI21_X1 _21140_ ( .A(_06133_ ), .B1(_02485_ ), .B2(_05731_ ), .ZN(_06134_ ) );
OAI22_X1 _21141_ ( .A1(_05916_ ), .A2(_06063_ ), .B1(_02484_ ), .B2(_06130_ ), .ZN(_06135_ ) );
AOI21_X1 _21142_ ( .A(_06134_ ), .B1(_06135_ ), .B2(_06102_ ), .ZN(_06136_ ) );
BUF_X4 _21143_ ( .A(_06074_ ), .Z(_06137_ ) );
NOR2_X1 _21144_ ( .A1(_06136_ ), .A2(_06137_ ), .ZN(_00021_ ) );
OAI22_X1 _21145_ ( .A1(_09806_ ), .A2(_05731_ ), .B1(_09105_ ), .B2(_09003_ ), .ZN(_06138_ ) );
OAI22_X1 _21146_ ( .A1(_05916_ ), .A2(_06063_ ), .B1(_09806_ ), .B2(_06130_ ), .ZN(_06139_ ) );
AOI21_X1 _21147_ ( .A(_06138_ ), .B1(_06139_ ), .B2(_06102_ ), .ZN(_06140_ ) );
NOR2_X1 _21148_ ( .A1(_06140_ ), .A2(_06137_ ), .ZN(_00022_ ) );
NAND2_X1 _21149_ ( .A1(_08908_ ), .A2(_09048_ ), .ZN(_06141_ ) );
OAI21_X1 _21150_ ( .A(_06141_ ), .B1(_09667_ ), .B2(_05731_ ), .ZN(_06142_ ) );
BUF_X4 _21151_ ( .A(_08995_ ), .Z(_06143_ ) );
BUF_X4 _21152_ ( .A(_09483_ ), .Z(_06144_ ) );
BUF_X4 _21153_ ( .A(_05808_ ), .Z(_06145_ ) );
CLKBUF_X2 _21154_ ( .A(_06018_ ), .Z(_06146_ ) );
NAND3_X1 _21155_ ( .A1(_06145_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06146_ ), .ZN(_06147_ ) );
INV_X1 _21156_ ( .A(_06147_ ), .ZN(_06148_ ) );
BUF_X4 _21157_ ( .A(_09122_ ), .Z(_06149_ ) );
BUF_X4 _21158_ ( .A(_09528_ ), .Z(_06150_ ) );
AOI221_X4 _21159_ ( .A(_06148_ ), .B1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06149_ ), .C1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06150_ ), .ZN(_06151_ ) );
BUF_X4 _21160_ ( .A(_09070_ ), .Z(_06152_ ) );
BUF_X4 _21161_ ( .A(_09093_ ), .Z(_06153_ ) );
BUF_X4 _21162_ ( .A(_06153_ ), .Z(_06154_ ) );
NAND3_X1 _21163_ ( .A1(_06152_ ), .A2(_06154_ ), .A3(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06155_ ) );
AOI21_X1 _21164_ ( .A(_06144_ ), .B1(_06151_ ), .B2(_06155_ ), .ZN(_06156_ ) );
BUF_X8 _21165_ ( .A(_05744_ ), .Z(_06157_ ) );
BUF_X4 _21166_ ( .A(_06157_ ), .Z(_06158_ ) );
BUF_X2 _21167_ ( .A(_09067_ ), .Z(_06159_ ) );
BUF_X4 _21168_ ( .A(_06018_ ), .Z(_06160_ ) );
NAND3_X1 _21169_ ( .A1(_06159_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06160_ ), .ZN(_06161_ ) );
INV_X1 _21170_ ( .A(_06161_ ), .ZN(_06162_ ) );
BUF_X4 _21171_ ( .A(_05865_ ), .Z(_06163_ ) );
AOI221_X4 _21172_ ( .A(_06162_ ), .B1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_09122_ ), .C1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06163_ ), .ZN(_06164_ ) );
BUF_X4 _21173_ ( .A(_09069_ ), .Z(_06165_ ) );
BUF_X4 _21174_ ( .A(_06165_ ), .Z(_06166_ ) );
BUF_X4 _21175_ ( .A(_06153_ ), .Z(_06167_ ) );
NAND3_X1 _21176_ ( .A1(_06166_ ), .A2(_06167_ ), .A3(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06168_ ) );
AOI21_X1 _21177_ ( .A(_06158_ ), .B1(_06164_ ), .B2(_06168_ ), .ZN(_06169_ ) );
NOR3_X1 _21178_ ( .A1(_06156_ ), .A2(_06169_ ), .A3(_09482_ ), .ZN(_06170_ ) );
NAND3_X1 _21179_ ( .A1(_06159_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06160_ ), .ZN(_06171_ ) );
INV_X1 _21180_ ( .A(_06171_ ), .ZN(_06172_ ) );
AOI221_X4 _21181_ ( .A(_06172_ ), .B1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_09122_ ), .C1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06163_ ), .ZN(_06173_ ) );
NAND3_X1 _21182_ ( .A1(_06166_ ), .A2(_06167_ ), .A3(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06174_ ) );
AOI21_X1 _21183_ ( .A(_06158_ ), .B1(_06173_ ), .B2(_06174_ ), .ZN(_06175_ ) );
BUF_X4 _21184_ ( .A(_09554_ ), .Z(_06176_ ) );
BUF_X4 _21185_ ( .A(_06176_ ), .Z(_06177_ ) );
BUF_X4 _21186_ ( .A(_09122_ ), .Z(_06178_ ) );
BUF_X4 _21187_ ( .A(_06178_ ), .Z(_06179_ ) );
AOI22_X1 _21188_ ( .A1(_06177_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06179_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06180_ ) );
BUF_X4 _21189_ ( .A(_09626_ ), .Z(_06181_ ) );
AOI22_X1 _21190_ ( .A1(_06181_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_09529_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06182_ ) );
AOI21_X1 _21191_ ( .A(_09084_ ), .B1(_06180_ ), .B2(_06182_ ), .ZN(_06183_ ) );
NOR3_X1 _21192_ ( .A1(_06175_ ), .A2(_09550_ ), .A3(_06183_ ), .ZN(_06184_ ) );
NOR3_X1 _21193_ ( .A1(_06170_ ), .A2(_06184_ ), .A3(_09665_ ), .ZN(_06185_ ) );
BUF_X4 _21194_ ( .A(_09046_ ), .Z(_06186_ ) );
CLKBUF_X2 _21195_ ( .A(_05765_ ), .Z(_06187_ ) );
AND3_X1 _21196_ ( .A1(_10429_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06187_ ), .ZN(_06188_ ) );
BUF_X4 _21197_ ( .A(_05865_ ), .Z(_06189_ ) );
BUF_X4 _21198_ ( .A(_09553_ ), .Z(_06190_ ) );
AOI221_X4 _21199_ ( .A(_06188_ ), .B1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06189_ ), .C1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06190_ ), .ZN(_06191_ ) );
BUF_X4 _21200_ ( .A(_09483_ ), .Z(_06192_ ) );
BUF_X4 _21201_ ( .A(_06165_ ), .Z(_06193_ ) );
BUF_X4 _21202_ ( .A(_06153_ ), .Z(_06194_ ) );
NAND3_X1 _21203_ ( .A1(_06193_ ), .A2(_06194_ ), .A3(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06195_ ) );
NAND3_X1 _21204_ ( .A1(_06191_ ), .A2(_06192_ ), .A3(_06195_ ), .ZN(_06196_ ) );
BUF_X4 _21205_ ( .A(_09119_ ), .Z(_06197_ ) );
BUF_X4 _21206_ ( .A(_06197_ ), .Z(_06198_ ) );
BUF_X4 _21207_ ( .A(_05809_ ), .Z(_06199_ ) );
MUX2_X1 _21208_ ( .A(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .S(_06199_ ), .Z(_06200_ ) );
MUX2_X1 _21209_ ( .A(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .S(_06199_ ), .Z(_06201_ ) );
MUX2_X1 _21210_ ( .A(_06200_ ), .B(_06201_ ), .S(_10431_ ), .Z(_06202_ ) );
OAI211_X1 _21211_ ( .A(_06196_ ), .B(_09463_ ), .C1(_06198_ ), .C2(_06202_ ), .ZN(_06203_ ) );
BUF_X4 _21212_ ( .A(_09481_ ), .Z(_06204_ ) );
BUF_X4 _21213_ ( .A(_09745_ ), .Z(_06205_ ) );
BUF_X4 _21214_ ( .A(_09626_ ), .Z(_06206_ ) );
BUF_X4 _21215_ ( .A(_06206_ ), .Z(_06207_ ) );
AOI22_X1 _21216_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06205_ ), .B1(_06207_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06208_ ) );
BUF_X4 _21217_ ( .A(_06157_ ), .Z(_06209_ ) );
BUF_X8 _21218_ ( .A(_09122_ ), .Z(_06210_ ) );
BUF_X4 _21219_ ( .A(_06210_ ), .Z(_06211_ ) );
BUF_X4 _21220_ ( .A(_09528_ ), .Z(_06212_ ) );
BUF_X4 _21221_ ( .A(_06212_ ), .Z(_06213_ ) );
AOI22_X1 _21222_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06211_ ), .B1(_06213_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06214_ ) );
NAND3_X1 _21223_ ( .A1(_06208_ ), .A2(_06209_ ), .A3(_06214_ ), .ZN(_06215_ ) );
BUF_X4 _21224_ ( .A(_09745_ ), .Z(_06216_ ) );
BUF_X4 _21225_ ( .A(_06206_ ), .Z(_06217_ ) );
AOI22_X1 _21226_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06216_ ), .B1(_06217_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06218_ ) );
BUF_X4 _21227_ ( .A(_09483_ ), .Z(_06219_ ) );
BUF_X4 _21228_ ( .A(_06210_ ), .Z(_06220_ ) );
BUF_X4 _21229_ ( .A(_06212_ ), .Z(_06221_ ) );
AOI22_X1 _21230_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06220_ ), .B1(_06221_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06222_ ) );
NAND3_X1 _21231_ ( .A1(_06218_ ), .A2(_06219_ ), .A3(_06222_ ), .ZN(_06223_ ) );
NAND3_X1 _21232_ ( .A1(_06204_ ), .A2(_06215_ ), .A3(_06223_ ), .ZN(_06224_ ) );
AOI21_X1 _21233_ ( .A(_06186_ ), .B1(_06203_ ), .B2(_06224_ ), .ZN(_06225_ ) );
OAI21_X1 _21234_ ( .A(_06143_ ), .B1(_06185_ ), .B2(_06225_ ), .ZN(_06226_ ) );
BUF_X4 _21235_ ( .A(_08993_ ), .Z(_06227_ ) );
CLKBUF_X2 _21236_ ( .A(_05748_ ), .Z(_06228_ ) );
BUF_X2 _21237_ ( .A(_06018_ ), .Z(_06229_ ) );
AND3_X1 _21238_ ( .A1(_06228_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06229_ ), .ZN(_06230_ ) );
BUF_X4 _21239_ ( .A(_05865_ ), .Z(_06231_ ) );
BUF_X4 _21240_ ( .A(_09554_ ), .Z(_06232_ ) );
AOI221_X4 _21241_ ( .A(_06230_ ), .B1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06231_ ), .C1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06232_ ), .ZN(_06233_ ) );
BUF_X2 _21242_ ( .A(_09483_ ), .Z(_06234_ ) );
BUF_X4 _21243_ ( .A(_09070_ ), .Z(_06235_ ) );
BUF_X4 _21244_ ( .A(_09094_ ), .Z(_06236_ ) );
NAND3_X1 _21245_ ( .A1(_06235_ ), .A2(_06236_ ), .A3(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06237_ ) );
NAND3_X1 _21246_ ( .A1(_06233_ ), .A2(_06234_ ), .A3(_06237_ ), .ZN(_06238_ ) );
BUF_X2 _21247_ ( .A(_05764_ ), .Z(_06239_ ) );
CLKBUF_X2 _21248_ ( .A(_06018_ ), .Z(_06240_ ) );
AND3_X1 _21249_ ( .A1(_06239_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06240_ ), .ZN(_06241_ ) );
BUF_X4 _21250_ ( .A(_05865_ ), .Z(_06242_ ) );
AOI221_X4 _21251_ ( .A(_06241_ ), .B1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06242_ ), .C1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C2(_09627_ ), .ZN(_06243_ ) );
BUF_X4 _21252_ ( .A(_05744_ ), .Z(_06244_ ) );
BUF_X4 _21253_ ( .A(_06244_ ), .Z(_06245_ ) );
BUF_X4 _21254_ ( .A(_10431_ ), .Z(_06246_ ) );
BUF_X4 _21255_ ( .A(_05809_ ), .Z(_06247_ ) );
BUF_X4 _21256_ ( .A(_06247_ ), .Z(_06248_ ) );
BUF_X4 _21257_ ( .A(_06248_ ), .Z(_06249_ ) );
NAND3_X1 _21258_ ( .A1(_06246_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06249_ ), .ZN(_06250_ ) );
NAND3_X1 _21259_ ( .A1(_06243_ ), .A2(_06245_ ), .A3(_06250_ ), .ZN(_06251_ ) );
BUF_X4 _21260_ ( .A(_09055_ ), .Z(_06252_ ) );
NAND3_X1 _21261_ ( .A1(_06238_ ), .A2(_06251_ ), .A3(_06252_ ), .ZN(_06253_ ) );
BUF_X4 _21262_ ( .A(_09481_ ), .Z(_06254_ ) );
BUF_X4 _21263_ ( .A(_09119_ ), .Z(_06255_ ) );
BUF_X2 _21264_ ( .A(_06018_ ), .Z(_06256_ ) );
NAND3_X1 _21265_ ( .A1(_06239_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06256_ ), .ZN(_06257_ ) );
INV_X1 _21266_ ( .A(_06257_ ), .ZN(_06258_ ) );
BUF_X4 _21267_ ( .A(_09528_ ), .Z(_06259_ ) );
AOI221_X4 _21268_ ( .A(_06258_ ), .B1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06178_ ), .C1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06259_ ), .ZN(_06260_ ) );
NAND3_X1 _21269_ ( .A1(_06193_ ), .A2(_06194_ ), .A3(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06261_ ) );
AOI21_X1 _21270_ ( .A(_06255_ ), .B1(_06260_ ), .B2(_06261_ ), .ZN(_06262_ ) );
BUF_X4 _21271_ ( .A(_06206_ ), .Z(_06263_ ) );
BUF_X4 _21272_ ( .A(_09123_ ), .Z(_06264_ ) );
AOI22_X1 _21273_ ( .A1(_06263_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06264_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06265_ ) );
BUF_X4 _21274_ ( .A(_09554_ ), .Z(_06266_ ) );
BUF_X4 _21275_ ( .A(_06266_ ), .Z(_06267_ ) );
BUF_X4 _21276_ ( .A(_06150_ ), .Z(_06268_ ) );
AOI22_X1 _21277_ ( .A1(_06267_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06268_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06269_ ) );
AOI21_X1 _21278_ ( .A(_06158_ ), .B1(_06265_ ), .B2(_06269_ ), .ZN(_06270_ ) );
OAI21_X1 _21279_ ( .A(_06254_ ), .B1(_06262_ ), .B2(_06270_ ), .ZN(_06271_ ) );
AOI21_X1 _21280_ ( .A(_09665_ ), .B1(_06253_ ), .B2(_06271_ ), .ZN(_06272_ ) );
AOI22_X1 _21281_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06205_ ), .B1(_06207_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06273_ ) );
BUF_X4 _21282_ ( .A(_06212_ ), .Z(_06274_ ) );
AOI22_X1 _21283_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06211_ ), .B1(_06274_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06275_ ) );
NAND3_X1 _21284_ ( .A1(_06273_ ), .A2(_06209_ ), .A3(_06275_ ), .ZN(_06276_ ) );
AOI22_X1 _21285_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06216_ ), .B1(_06217_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06277_ ) );
AOI22_X1 _21286_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06220_ ), .B1(_06221_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06278_ ) );
NAND3_X1 _21287_ ( .A1(_06277_ ), .A2(_06219_ ), .A3(_06278_ ), .ZN(_06279_ ) );
NAND3_X1 _21288_ ( .A1(_06204_ ), .A2(_06276_ ), .A3(_06279_ ), .ZN(_06280_ ) );
AOI22_X1 _21289_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06267_ ), .B1(_09795_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06281_ ) );
AOI22_X1 _21290_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_09484_ ), .B1(_06268_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06282_ ) );
AOI21_X1 _21291_ ( .A(_06197_ ), .B1(_06281_ ), .B2(_06282_ ), .ZN(_06283_ ) );
BUF_X4 _21292_ ( .A(_05744_ ), .Z(_06284_ ) );
BUF_X4 _21293_ ( .A(_09554_ ), .Z(_06285_ ) );
BUF_X4 _21294_ ( .A(_06285_ ), .Z(_06286_ ) );
AOI22_X1 _21295_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06286_ ), .B1(_06181_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06287_ ) );
BUF_X4 _21296_ ( .A(_09123_ ), .Z(_06288_ ) );
BUF_X4 _21297_ ( .A(_06163_ ), .Z(_06289_ ) );
AOI22_X1 _21298_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06288_ ), .B1(_06289_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06290_ ) );
AOI21_X1 _21299_ ( .A(_06284_ ), .B1(_06287_ ), .B2(_06290_ ), .ZN(_06291_ ) );
OAI21_X1 _21300_ ( .A(_09463_ ), .B1(_06283_ ), .B2(_06291_ ), .ZN(_06292_ ) );
AOI21_X1 _21301_ ( .A(_06186_ ), .B1(_06280_ ), .B2(_06292_ ), .ZN(_06293_ ) );
OAI21_X1 _21302_ ( .A(_06227_ ), .B1(_06272_ ), .B2(_06293_ ), .ZN(_06294_ ) );
AOI21_X1 _21303_ ( .A(_02457_ ), .B1(_06226_ ), .B2(_06294_ ), .ZN(_06295_ ) );
BUF_X2 _21304_ ( .A(_05766_ ), .Z(_06296_ ) );
AND3_X1 _21305_ ( .A1(_10430_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06296_ ), .ZN(_06297_ ) );
BUF_X4 _21306_ ( .A(_09554_ ), .Z(_06298_ ) );
AOI221_X4 _21307_ ( .A(_06297_ ), .B1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06163_ ), .C1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06298_ ), .ZN(_06299_ ) );
BUF_X4 _21308_ ( .A(_06244_ ), .Z(_06300_ ) );
NAND3_X1 _21309_ ( .A1(_09071_ ), .A2(_09095_ ), .A3(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06301_ ) );
NAND3_X1 _21310_ ( .A1(_06299_ ), .A2(_06300_ ), .A3(_06301_ ), .ZN(_06302_ ) );
BUF_X4 _21311_ ( .A(_09055_ ), .Z(_06303_ ) );
BUF_X4 _21312_ ( .A(_09554_ ), .Z(_06304_ ) );
BUF_X4 _21313_ ( .A(_06304_ ), .Z(_06305_ ) );
BUF_X4 _21314_ ( .A(_09529_ ), .Z(_06306_ ) );
AOI22_X1 _21315_ ( .A1(_06305_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06306_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06307_ ) );
BUF_X4 _21316_ ( .A(_09084_ ), .Z(_06308_ ) );
BUF_X4 _21317_ ( .A(_09070_ ), .Z(_06309_ ) );
NAND3_X1 _21318_ ( .A1(_06309_ ), .A2(_06154_ ), .A3(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06310_ ) );
BUF_X4 _21319_ ( .A(_06248_ ), .Z(_06311_ ) );
NAND3_X1 _21320_ ( .A1(_06246_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06311_ ), .ZN(_06312_ ) );
NAND4_X1 _21321_ ( .A1(_06307_ ), .A2(_06308_ ), .A3(_06310_ ), .A4(_06312_ ), .ZN(_06313_ ) );
NAND3_X1 _21322_ ( .A1(_06302_ ), .A2(_06303_ ), .A3(_06313_ ), .ZN(_06314_ ) );
BUF_X4 _21323_ ( .A(_09481_ ), .Z(_06315_ ) );
BUF_X4 _21324_ ( .A(_06304_ ), .Z(_06316_ ) );
BUF_X4 _21325_ ( .A(_09626_ ), .Z(_06317_ ) );
BUF_X4 _21326_ ( .A(_06317_ ), .Z(_06318_ ) );
AOI22_X1 _21327_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06316_ ), .B1(_06318_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06319_ ) );
BUF_X4 _21328_ ( .A(_06244_ ), .Z(_06320_ ) );
BUF_X4 _21329_ ( .A(_06210_ ), .Z(_06321_ ) );
BUF_X4 _21330_ ( .A(_09529_ ), .Z(_06322_ ) );
AOI22_X1 _21331_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06321_ ), .B1(_06322_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06323_ ) );
NAND3_X1 _21332_ ( .A1(_06319_ ), .A2(_06320_ ), .A3(_06323_ ), .ZN(_06324_ ) );
BUF_X4 _21333_ ( .A(_06210_ ), .Z(_06325_ ) );
BUF_X4 _21334_ ( .A(_09528_ ), .Z(_06326_ ) );
BUF_X4 _21335_ ( .A(_06326_ ), .Z(_06327_ ) );
AOI22_X1 _21336_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06325_ ), .B1(_06327_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06328_ ) );
BUF_X4 _21337_ ( .A(_09483_ ), .Z(_06329_ ) );
BUF_X4 _21338_ ( .A(_06165_ ), .Z(_06330_ ) );
BUF_X4 _21339_ ( .A(_06153_ ), .Z(_06331_ ) );
NAND3_X1 _21340_ ( .A1(_06330_ ), .A2(_06331_ ), .A3(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06332_ ) );
BUF_X4 _21341_ ( .A(_06248_ ), .Z(_06333_ ) );
NAND3_X1 _21342_ ( .A1(_06193_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06333_ ), .ZN(_06334_ ) );
NAND4_X1 _21343_ ( .A1(_06328_ ), .A2(_06329_ ), .A3(_06332_ ), .A4(_06334_ ), .ZN(_06335_ ) );
NAND3_X1 _21344_ ( .A1(_06315_ ), .A2(_06324_ ), .A3(_06335_ ), .ZN(_06336_ ) );
NAND3_X1 _21345_ ( .A1(_06314_ ), .A2(_11056_ ), .A3(_06336_ ), .ZN(_06337_ ) );
BUF_X4 _21346_ ( .A(_08995_ ), .Z(_06338_ ) );
BUF_X4 _21347_ ( .A(_06179_ ), .Z(_06339_ ) );
BUF_X4 _21348_ ( .A(_09529_ ), .Z(_06340_ ) );
AOI22_X1 _21349_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06339_ ), .B1(_06340_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06341_ ) );
BUF_X4 _21350_ ( .A(_09745_ ), .Z(_06342_ ) );
BUF_X4 _21351_ ( .A(_06206_ ), .Z(_06343_ ) );
AOI22_X1 _21352_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06342_ ), .B1(_06343_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06344_ ) );
NAND3_X1 _21353_ ( .A1(_06341_ ), .A2(_06320_ ), .A3(_06344_ ), .ZN(_06345_ ) );
BUF_X4 _21354_ ( .A(_09745_ ), .Z(_06346_ ) );
BUF_X4 _21355_ ( .A(_06210_ ), .Z(_06347_ ) );
AOI22_X1 _21356_ ( .A1(_06346_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06347_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06348_ ) );
NAND3_X1 _21357_ ( .A1(_06330_ ), .A2(_06331_ ), .A3(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06349_ ) );
BUF_X4 _21358_ ( .A(_06153_ ), .Z(_06350_ ) );
BUF_X4 _21359_ ( .A(_05868_ ), .Z(_06351_ ) );
BUF_X4 _21360_ ( .A(_06351_ ), .Z(_06352_ ) );
BUF_X4 _21361_ ( .A(_06352_ ), .Z(_06353_ ) );
BUF_X4 _21362_ ( .A(_05869_ ), .Z(_06354_ ) );
BUF_X4 _21363_ ( .A(_06354_ ), .Z(_06355_ ) );
BUF_X4 _21364_ ( .A(_06355_ ), .Z(_06356_ ) );
OAI211_X1 _21365_ ( .A(_06350_ ), .B(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06353_ ), .C2(_06356_ ), .ZN(_06357_ ) );
NAND4_X1 _21366_ ( .A1(_06348_ ), .A2(_06329_ ), .A3(_06349_ ), .A4(_06357_ ), .ZN(_06358_ ) );
NAND3_X1 _21367_ ( .A1(_06315_ ), .A2(_06345_ ), .A3(_06358_ ), .ZN(_06359_ ) );
BUF_X4 _21368_ ( .A(_09529_ ), .Z(_06360_ ) );
AOI22_X1 _21369_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06321_ ), .B1(_06360_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06361_ ) );
BUF_X4 _21370_ ( .A(_09483_ ), .Z(_06362_ ) );
AOI22_X1 _21371_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06216_ ), .B1(_06217_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06363_ ) );
NAND3_X1 _21372_ ( .A1(_06361_ ), .A2(_06362_ ), .A3(_06363_ ), .ZN(_06364_ ) );
BUF_X4 _21373_ ( .A(_09745_ ), .Z(_06365_ ) );
BUF_X4 _21374_ ( .A(_06206_ ), .Z(_06366_ ) );
AOI22_X1 _21375_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06365_ ), .B1(_06366_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06367_ ) );
BUF_X4 _21376_ ( .A(_06244_ ), .Z(_06368_ ) );
BUF_X4 _21377_ ( .A(_06210_ ), .Z(_06369_ ) );
BUF_X4 _21378_ ( .A(_06326_ ), .Z(_06370_ ) );
AOI22_X1 _21379_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06369_ ), .B1(_06370_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06371_ ) );
NAND3_X1 _21380_ ( .A1(_06367_ ), .A2(_06368_ ), .A3(_06371_ ), .ZN(_06372_ ) );
NAND3_X1 _21381_ ( .A1(_09056_ ), .A2(_06364_ ), .A3(_06372_ ), .ZN(_06373_ ) );
NAND3_X1 _21382_ ( .A1(_06359_ ), .A2(_09487_ ), .A3(_06373_ ), .ZN(_06374_ ) );
NAND3_X1 _21383_ ( .A1(_06337_ ), .A2(_06338_ ), .A3(_06374_ ), .ZN(_06375_ ) );
AOI22_X1 _21384_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06205_ ), .B1(_06207_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06376_ ) );
AOI22_X1 _21385_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06211_ ), .B1(_06213_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06377_ ) );
NAND3_X1 _21386_ ( .A1(_06376_ ), .A2(_06209_ ), .A3(_06377_ ), .ZN(_06378_ ) );
BUF_X4 _21387_ ( .A(_06210_ ), .Z(_06379_ ) );
BUF_X4 _21388_ ( .A(_06326_ ), .Z(_06380_ ) );
AOI22_X1 _21389_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06379_ ), .B1(_06380_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06381_ ) );
BUF_X4 _21390_ ( .A(_06298_ ), .Z(_06382_ ) );
BUF_X4 _21391_ ( .A(_09626_ ), .Z(_06383_ ) );
BUF_X4 _21392_ ( .A(_06383_ ), .Z(_06384_ ) );
AOI22_X1 _21393_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06382_ ), .B1(_06384_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06385_ ) );
NAND3_X1 _21394_ ( .A1(_06381_ ), .A2(_06219_ ), .A3(_06385_ ), .ZN(_06386_ ) );
NAND3_X1 _21395_ ( .A1(_06204_ ), .A2(_06378_ ), .A3(_06386_ ), .ZN(_06387_ ) );
BUF_X4 _21396_ ( .A(_09055_ ), .Z(_06388_ ) );
AOI22_X1 _21397_ ( .A1(_06263_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06264_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06389_ ) );
BUF_X4 _21398_ ( .A(_06157_ ), .Z(_06390_ ) );
CLKBUF_X2 _21399_ ( .A(_09091_ ), .Z(_06391_ ) );
BUF_X2 _21400_ ( .A(_06391_ ), .Z(_06392_ ) );
BUF_X4 _21401_ ( .A(_06392_ ), .Z(_06393_ ) );
BUF_X4 _21402_ ( .A(_06352_ ), .Z(_06394_ ) );
BUF_X4 _21403_ ( .A(_06354_ ), .Z(_06395_ ) );
OAI211_X1 _21404_ ( .A(_06393_ ), .B(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06394_ ), .C2(_06395_ ), .ZN(_06396_ ) );
BUF_X4 _21405_ ( .A(_09069_ ), .Z(_06397_ ) );
BUF_X4 _21406_ ( .A(_06397_ ), .Z(_06398_ ) );
BUF_X4 _21407_ ( .A(_05809_ ), .Z(_06399_ ) );
BUF_X4 _21408_ ( .A(_06399_ ), .Z(_06400_ ) );
BUF_X4 _21409_ ( .A(_06400_ ), .Z(_06401_ ) );
NAND3_X1 _21410_ ( .A1(_06398_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06401_ ), .ZN(_06402_ ) );
NAND4_X1 _21411_ ( .A1(_06389_ ), .A2(_06390_ ), .A3(_06396_ ), .A4(_06402_ ), .ZN(_06403_ ) );
AOI22_X1 _21412_ ( .A1(_06207_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06264_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06404_ ) );
BUF_X4 _21413_ ( .A(_09119_ ), .Z(_06405_ ) );
OAI211_X1 _21414_ ( .A(_06393_ ), .B(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06394_ ), .C2(_06395_ ), .ZN(_06406_ ) );
BUF_X4 _21415_ ( .A(_06397_ ), .Z(_06407_ ) );
BUF_X4 _21416_ ( .A(_06400_ ), .Z(_06408_ ) );
NAND3_X1 _21417_ ( .A1(_06407_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06408_ ), .ZN(_06409_ ) );
NAND4_X1 _21418_ ( .A1(_06404_ ), .A2(_06405_ ), .A3(_06406_ ), .A4(_06409_ ), .ZN(_06410_ ) );
NAND3_X1 _21419_ ( .A1(_06388_ ), .A2(_06403_ ), .A3(_06410_ ), .ZN(_06411_ ) );
AOI21_X1 _21420_ ( .A(_06186_ ), .B1(_06387_ ), .B2(_06411_ ), .ZN(_06412_ ) );
BUF_X4 _21421_ ( .A(_09664_ ), .Z(_06413_ ) );
BUF_X4 _21422_ ( .A(_09481_ ), .Z(_06414_ ) );
AOI22_X1 _21423_ ( .A1(_06207_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06288_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06415_ ) );
NAND3_X1 _21424_ ( .A1(_06407_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06401_ ), .ZN(_06416_ ) );
BUF_X4 _21425_ ( .A(_06351_ ), .Z(_06417_ ) );
BUF_X4 _21426_ ( .A(_06354_ ), .Z(_06418_ ) );
OAI211_X1 _21427_ ( .A(_06393_ ), .B(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06417_ ), .C2(_06418_ ), .ZN(_06419_ ) );
NAND4_X1 _21428_ ( .A1(_06415_ ), .A2(_06390_ ), .A3(_06416_ ), .A4(_06419_ ), .ZN(_06420_ ) );
BUF_X4 _21429_ ( .A(_09745_ ), .Z(_06421_ ) );
BUF_X4 _21430_ ( .A(_09123_ ), .Z(_06422_ ) );
AOI22_X1 _21431_ ( .A1(_06421_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06422_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06423_ ) );
BUF_X4 _21432_ ( .A(_09528_ ), .Z(_06424_ ) );
BUF_X4 _21433_ ( .A(_06424_ ), .Z(_06425_ ) );
AOI22_X1 _21434_ ( .A1(_06366_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06425_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06426_ ) );
NAND3_X1 _21435_ ( .A1(_06423_ ), .A2(_06426_ ), .A3(_06255_ ), .ZN(_06427_ ) );
NAND3_X1 _21436_ ( .A1(_06414_ ), .A2(_06420_ ), .A3(_06427_ ), .ZN(_06428_ ) );
BUF_X4 _21437_ ( .A(_06383_ ), .Z(_06429_ ) );
BUF_X4 _21438_ ( .A(_09122_ ), .Z(_06430_ ) );
BUF_X4 _21439_ ( .A(_06430_ ), .Z(_06431_ ) );
AOI22_X1 _21440_ ( .A1(_06429_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06431_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06432_ ) );
BUF_X4 _21441_ ( .A(_06157_ ), .Z(_06433_ ) );
BUF_X2 _21442_ ( .A(_06145_ ), .Z(_06434_ ) );
BUF_X4 _21443_ ( .A(_06434_ ), .Z(_06435_ ) );
BUF_X2 _21444_ ( .A(_06296_ ), .Z(_06436_ ) );
BUF_X4 _21445_ ( .A(_06436_ ), .Z(_06437_ ) );
NAND3_X1 _21446_ ( .A1(_06435_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06437_ ), .ZN(_06438_ ) );
CLKBUF_X2 _21447_ ( .A(_05748_ ), .Z(_06439_ ) );
BUF_X2 _21448_ ( .A(_06439_ ), .Z(_06440_ ) );
BUF_X4 _21449_ ( .A(_06440_ ), .Z(_06441_ ) );
NAND3_X1 _21450_ ( .A1(_06441_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06393_ ), .ZN(_06442_ ) );
NAND4_X1 _21451_ ( .A1(_06432_ ), .A2(_06433_ ), .A3(_06438_ ), .A4(_06442_ ), .ZN(_06443_ ) );
BUF_X4 _21452_ ( .A(_06232_ ), .Z(_06444_ ) );
BUF_X4 _21453_ ( .A(_06259_ ), .Z(_06445_ ) );
AOI22_X1 _21454_ ( .A1(_06444_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06445_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06446_ ) );
NAND3_X1 _21455_ ( .A1(_06435_ ), .A2(_06393_ ), .A3(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06447_ ) );
BUF_X4 _21456_ ( .A(_10430_ ), .Z(_06448_ ) );
NAND3_X1 _21457_ ( .A1(_06448_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06437_ ), .ZN(_06449_ ) );
NAND4_X1 _21458_ ( .A1(_06446_ ), .A2(_06197_ ), .A3(_06447_ ), .A4(_06449_ ), .ZN(_06450_ ) );
NAND3_X1 _21459_ ( .A1(_09463_ ), .A2(_06443_ ), .A3(_06450_ ), .ZN(_06451_ ) );
AOI21_X1 _21460_ ( .A(_06413_ ), .B1(_06428_ ), .B2(_06451_ ), .ZN(_06452_ ) );
OAI21_X1 _21461_ ( .A(_06227_ ), .B1(_06412_ ), .B2(_06452_ ), .ZN(_06453_ ) );
AOI21_X1 _21462_ ( .A(_09604_ ), .B1(_06375_ ), .B2(_06453_ ), .ZN(_06454_ ) );
OAI21_X1 _21463_ ( .A(_09493_ ), .B1(_06295_ ), .B2(_06454_ ), .ZN(_06455_ ) );
CLKBUF_X2 _21464_ ( .A(_05748_ ), .Z(_06456_ ) );
AND3_X1 _21465_ ( .A1(_06456_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06187_ ), .ZN(_06457_ ) );
AOI221_X4 _21466_ ( .A(_06457_ ), .B1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06189_ ), .C1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06190_ ), .ZN(_06458_ ) );
BUF_X4 _21467_ ( .A(_06165_ ), .Z(_06459_ ) );
BUF_X4 _21468_ ( .A(_06153_ ), .Z(_06460_ ) );
NAND3_X1 _21469_ ( .A1(_06459_ ), .A2(_06460_ ), .A3(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06461_ ) );
NAND3_X1 _21470_ ( .A1(_06458_ ), .A2(_06329_ ), .A3(_06461_ ), .ZN(_06462_ ) );
BUF_X4 _21471_ ( .A(_09481_ ), .Z(_06463_ ) );
BUF_X4 _21472_ ( .A(_06160_ ), .Z(_06464_ ) );
MUX2_X1 _21473_ ( .A(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .S(_06464_ ), .Z(_06465_ ) );
MUX2_X1 _21474_ ( .A(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .S(_06464_ ), .Z(_06466_ ) );
MUX2_X1 _21475_ ( .A(_06465_ ), .B(_06466_ ), .S(_06448_ ), .Z(_06467_ ) );
OAI211_X1 _21476_ ( .A(_06462_ ), .B(_06463_ ), .C1(_06198_ ), .C2(_06467_ ), .ZN(_06468_ ) );
BUF_X4 _21477_ ( .A(_06317_ ), .Z(_06469_ ) );
BUF_X4 _21478_ ( .A(_09123_ ), .Z(_06470_ ) );
AOI22_X1 _21479_ ( .A1(_06469_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06470_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06471_ ) );
OAI211_X1 _21480_ ( .A(_06350_ ), .B(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06353_ ), .C2(_06356_ ), .ZN(_06472_ ) );
BUF_X4 _21481_ ( .A(_06165_ ), .Z(_06473_ ) );
NAND3_X1 _21482_ ( .A1(_06473_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06333_ ), .ZN(_06474_ ) );
NAND4_X1 _21483_ ( .A1(_06471_ ), .A2(_06192_ ), .A3(_06472_ ), .A4(_06474_ ), .ZN(_06475_ ) );
BUF_X4 _21484_ ( .A(_06317_ ), .Z(_06476_ ) );
BUF_X4 _21485_ ( .A(_09123_ ), .Z(_06477_ ) );
AOI22_X1 _21486_ ( .A1(_06476_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06477_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06478_ ) );
BUF_X2 _21487_ ( .A(_06157_ ), .Z(_06479_ ) );
BUF_X4 _21488_ ( .A(_06352_ ), .Z(_06480_ ) );
BUF_X4 _21489_ ( .A(_06355_ ), .Z(_06481_ ) );
OAI211_X1 _21490_ ( .A(_06350_ ), .B(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06480_ ), .C2(_06481_ ), .ZN(_06482_ ) );
BUF_X2 _21491_ ( .A(_06397_ ), .Z(_06483_ ) );
BUF_X2 _21492_ ( .A(_06400_ ), .Z(_06484_ ) );
NAND3_X1 _21493_ ( .A1(_06483_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06484_ ), .ZN(_06485_ ) );
NAND4_X1 _21494_ ( .A1(_06478_ ), .A2(_06479_ ), .A3(_06482_ ), .A4(_06485_ ), .ZN(_06486_ ) );
NAND3_X1 _21495_ ( .A1(_10050_ ), .A2(_06475_ ), .A3(_06486_ ), .ZN(_06487_ ) );
AOI21_X1 _21496_ ( .A(_09594_ ), .B1(_06468_ ), .B2(_06487_ ), .ZN(_06488_ ) );
OAI211_X1 _21497_ ( .A(_05809_ ), .B(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(_05868_ ), .C2(_05869_ ), .ZN(_06489_ ) );
INV_X1 _21498_ ( .A(_06489_ ), .ZN(_06490_ ) );
AOI221_X4 _21499_ ( .A(_06490_ ), .B1(_06189_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_09554_ ), .ZN(_06491_ ) );
BUF_X4 _21500_ ( .A(_06165_ ), .Z(_06492_ ) );
NAND3_X1 _21501_ ( .A1(_06492_ ), .A2(_06167_ ), .A3(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06493_ ) );
AOI21_X1 _21502_ ( .A(_06433_ ), .B1(_06491_ ), .B2(_06493_ ), .ZN(_06494_ ) );
BUF_X4 _21503_ ( .A(_09119_ ), .Z(_06495_ ) );
AOI22_X1 _21504_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06177_ ), .B1(_06181_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06496_ ) );
AOI22_X1 _21505_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06288_ ), .B1(_06289_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06497_ ) );
AOI21_X1 _21506_ ( .A(_06495_ ), .B1(_06496_ ), .B2(_06497_ ), .ZN(_06498_ ) );
OAI21_X1 _21507_ ( .A(_09482_ ), .B1(_06494_ ), .B2(_06498_ ), .ZN(_06499_ ) );
BUF_X4 _21508_ ( .A(_09055_ ), .Z(_06500_ ) );
AOI22_X1 _21509_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06286_ ), .B1(_06181_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06501_ ) );
AOI22_X1 _21510_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06264_ ), .B1(_06289_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06502_ ) );
AOI21_X1 _21511_ ( .A(_06495_ ), .B1(_06501_ ), .B2(_06502_ ), .ZN(_06503_ ) );
BUF_X4 _21512_ ( .A(_09626_ ), .Z(_06504_ ) );
AOI22_X1 _21513_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06304_ ), .B1(_06504_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06505_ ) );
BUF_X4 _21514_ ( .A(_06163_ ), .Z(_06506_ ) );
AOI22_X1 _21515_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06431_ ), .B1(_06506_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06507_ ) );
AOI21_X1 _21516_ ( .A(_06244_ ), .B1(_06505_ ), .B2(_06507_ ), .ZN(_06508_ ) );
OAI21_X1 _21517_ ( .A(_06500_ ), .B1(_06503_ ), .B2(_06508_ ), .ZN(_06509_ ) );
AOI21_X1 _21518_ ( .A(_06413_ ), .B1(_06499_ ), .B2(_06509_ ), .ZN(_06510_ ) );
NOR3_X1 _21519_ ( .A1(_06488_ ), .A2(_06227_ ), .A3(_06510_ ), .ZN(_06511_ ) );
AND3_X1 _21520_ ( .A1(_10429_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_05809_ ), .ZN(_06512_ ) );
AOI221_X4 _21521_ ( .A(_06512_ ), .B1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06189_ ), .C1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06190_ ), .ZN(_06513_ ) );
BUF_X4 _21522_ ( .A(_09483_ ), .Z(_06514_ ) );
BUF_X4 _21523_ ( .A(_06153_ ), .Z(_06515_ ) );
NAND3_X1 _21524_ ( .A1(_06473_ ), .A2(_06515_ ), .A3(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06516_ ) );
NAND3_X1 _21525_ ( .A1(_06513_ ), .A2(_06514_ ), .A3(_06516_ ), .ZN(_06517_ ) );
MUX2_X1 _21526_ ( .A(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .S(_06199_ ), .Z(_06518_ ) );
MUX2_X1 _21527_ ( .A(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .S(_06199_ ), .Z(_06519_ ) );
MUX2_X1 _21528_ ( .A(_06518_ ), .B(_06519_ ), .S(_10431_ ), .Z(_06520_ ) );
OAI211_X1 _21529_ ( .A(_06517_ ), .B(_09463_ ), .C1(_06198_ ), .C2(_06520_ ), .ZN(_06521_ ) );
BUF_X4 _21530_ ( .A(_06298_ ), .Z(_06522_ ) );
AOI22_X1 _21531_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06522_ ), .B1(_06384_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06523_ ) );
BUF_X4 _21532_ ( .A(_06424_ ), .Z(_06524_ ) );
AOI22_X1 _21533_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06477_ ), .B1(_06524_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06525_ ) );
AOI21_X1 _21534_ ( .A(_06390_ ), .B1(_06523_ ), .B2(_06525_ ), .ZN(_06526_ ) );
BUF_X4 _21535_ ( .A(_09627_ ), .Z(_06527_ ) );
AOI22_X1 _21536_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06444_ ), .B1(_06527_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06528_ ) );
AOI22_X1 _21537_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06422_ ), .B1(_06445_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06529_ ) );
AOI21_X1 _21538_ ( .A(_06197_ ), .B1(_06528_ ), .B2(_06529_ ), .ZN(_06530_ ) );
OAI21_X1 _21539_ ( .A(_06463_ ), .B1(_06526_ ), .B2(_06530_ ), .ZN(_06531_ ) );
AOI21_X1 _21540_ ( .A(_06413_ ), .B1(_06521_ ), .B2(_06531_ ), .ZN(_06532_ ) );
AOI22_X1 _21541_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06444_ ), .B1(_06527_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06533_ ) );
AOI22_X1 _21542_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06422_ ), .B1(_06445_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06534_ ) );
AOI21_X1 _21543_ ( .A(_06197_ ), .B1(_06533_ ), .B2(_06534_ ), .ZN(_06535_ ) );
AOI22_X1 _21544_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06177_ ), .B1(_06504_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06536_ ) );
AOI22_X1 _21545_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06431_ ), .B1(_06506_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06537_ ) );
AOI21_X1 _21546_ ( .A(_06284_ ), .B1(_06536_ ), .B2(_06537_ ), .ZN(_06538_ ) );
OAI21_X1 _21547_ ( .A(_09482_ ), .B1(_06535_ ), .B2(_06538_ ), .ZN(_06539_ ) );
BUF_X4 _21548_ ( .A(_06383_ ), .Z(_06540_ ) );
AOI22_X1 _21549_ ( .A1(_06540_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06431_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06541_ ) );
OAI211_X1 _21550_ ( .A(_09094_ ), .B(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06417_ ), .C2(_06418_ ), .ZN(_06542_ ) );
BUF_X4 _21551_ ( .A(_06296_ ), .Z(_06543_ ) );
BUF_X4 _21552_ ( .A(_06543_ ), .Z(_06544_ ) );
NAND3_X1 _21553_ ( .A1(_06435_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06544_ ), .ZN(_06545_ ) );
NAND4_X1 _21554_ ( .A1(_06541_ ), .A2(_06433_ ), .A3(_06542_ ), .A4(_06545_ ), .ZN(_06546_ ) );
AOI22_X1 _21555_ ( .A1(_06384_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06179_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06547_ ) );
OAI211_X1 _21556_ ( .A(_09094_ ), .B(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06417_ ), .C2(_06418_ ), .ZN(_06548_ ) );
NAND3_X1 _21557_ ( .A1(_06435_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06544_ ), .ZN(_06549_ ) );
NAND4_X1 _21558_ ( .A1(_06547_ ), .A2(_06495_ ), .A3(_06548_ ), .A4(_06549_ ), .ZN(_06550_ ) );
NAND3_X1 _21559_ ( .A1(_06500_ ), .A2(_06546_ ), .A3(_06550_ ), .ZN(_06551_ ) );
AOI21_X1 _21560_ ( .A(_10252_ ), .B1(_06539_ ), .B2(_06551_ ), .ZN(_06552_ ) );
NOR3_X1 _21561_ ( .A1(_06532_ ), .A2(_06552_ ), .A3(_08995_ ), .ZN(_06553_ ) );
OAI21_X1 _21562_ ( .A(_02409_ ), .B1(_06511_ ), .B2(_06553_ ), .ZN(_06554_ ) );
BUF_X4 _21563_ ( .A(_09055_ ), .Z(_06555_ ) );
BUF_X4 _21564_ ( .A(_09084_ ), .Z(_06556_ ) );
CLKBUF_X2 _21565_ ( .A(_05748_ ), .Z(_06557_ ) );
AND3_X1 _21566_ ( .A1(_06557_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06146_ ), .ZN(_06558_ ) );
BUF_X4 _21567_ ( .A(_05865_ ), .Z(_06559_ ) );
AOI221_X4 _21568_ ( .A(_06558_ ), .B1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06559_ ), .C1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06266_ ), .ZN(_06560_ ) );
BUF_X4 _21569_ ( .A(_09070_ ), .Z(_06561_ ) );
BUF_X4 _21570_ ( .A(_09094_ ), .Z(_06562_ ) );
NAND3_X1 _21571_ ( .A1(_06561_ ), .A2(_06562_ ), .A3(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06563_ ) );
AOI21_X1 _21572_ ( .A(_06556_ ), .B1(_06560_ ), .B2(_06563_ ), .ZN(_06564_ ) );
BUF_X4 _21573_ ( .A(_06157_ ), .Z(_06565_ ) );
AND3_X1 _21574_ ( .A1(_06228_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06256_ ), .ZN(_06566_ ) );
AOI221_X4 _21575_ ( .A(_06566_ ), .B1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06242_ ), .C1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06285_ ), .ZN(_06567_ ) );
BUF_X4 _21576_ ( .A(_09070_ ), .Z(_06568_ ) );
BUF_X4 _21577_ ( .A(_09094_ ), .Z(_06569_ ) );
NAND3_X1 _21578_ ( .A1(_06568_ ), .A2(_06569_ ), .A3(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06570_ ) );
AOI21_X1 _21579_ ( .A(_06565_ ), .B1(_06567_ ), .B2(_06570_ ), .ZN(_06571_ ) );
OAI21_X1 _21580_ ( .A(_06555_ ), .B1(_06564_ ), .B2(_06571_ ), .ZN(_06572_ ) );
BUF_X4 _21581_ ( .A(_09481_ ), .Z(_06573_ ) );
BUF_X4 _21582_ ( .A(_06304_ ), .Z(_06574_ ) );
AOI22_X1 _21583_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06574_ ), .B1(_06469_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06575_ ) );
BUF_X4 _21584_ ( .A(_09084_ ), .Z(_06576_ ) );
AOI22_X1 _21585_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06339_ ), .B1(_06340_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06577_ ) );
NAND3_X1 _21586_ ( .A1(_06575_ ), .A2(_06576_ ), .A3(_06577_ ), .ZN(_06578_ ) );
AOI22_X1 _21587_ ( .A1(_06574_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06321_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06579_ ) );
BUF_X4 _21588_ ( .A(_06504_ ), .Z(_06580_ ) );
AOI22_X1 _21589_ ( .A1(_06580_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06340_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06581_ ) );
BUF_X4 _21590_ ( .A(_06244_ ), .Z(_06582_ ) );
NAND3_X1 _21591_ ( .A1(_06579_ ), .A2(_06581_ ), .A3(_06582_ ), .ZN(_06583_ ) );
NAND3_X1 _21592_ ( .A1(_06573_ ), .A2(_06578_ ), .A3(_06583_ ), .ZN(_06584_ ) );
NAND3_X1 _21593_ ( .A1(_06572_ ), .A2(_09784_ ), .A3(_06584_ ), .ZN(_06585_ ) );
AOI22_X1 _21594_ ( .A1(_06580_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06379_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06586_ ) );
BUF_X4 _21595_ ( .A(_06352_ ), .Z(_06587_ ) );
BUF_X4 _21596_ ( .A(_06355_ ), .Z(_06588_ ) );
OAI211_X1 _21597_ ( .A(_06194_ ), .B(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06587_ ), .C2(_06588_ ), .ZN(_06589_ ) );
BUF_X4 _21598_ ( .A(_06248_ ), .Z(_06590_ ) );
NAND3_X1 _21599_ ( .A1(_06309_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06590_ ), .ZN(_06591_ ) );
NAND4_X1 _21600_ ( .A1(_06586_ ), .A2(_06556_ ), .A3(_06589_ ), .A4(_06591_ ), .ZN(_06592_ ) );
BUF_X4 _21601_ ( .A(_06317_ ), .Z(_06593_ ) );
BUF_X4 _21602_ ( .A(_06210_ ), .Z(_06594_ ) );
AOI22_X1 _21603_ ( .A1(_06593_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06594_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06595_ ) );
BUF_X4 _21604_ ( .A(_06244_ ), .Z(_06596_ ) );
NAND3_X1 _21605_ ( .A1(_06309_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06590_ ), .ZN(_06597_ ) );
BUF_X4 _21606_ ( .A(_09093_ ), .Z(_06598_ ) );
BUF_X2 _21607_ ( .A(_06598_ ), .Z(_06599_ ) );
BUF_X4 _21608_ ( .A(_06352_ ), .Z(_06600_ ) );
BUF_X4 _21609_ ( .A(_06355_ ), .Z(_06601_ ) );
OAI211_X1 _21610_ ( .A(_06599_ ), .B(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06600_ ), .C2(_06601_ ), .ZN(_06602_ ) );
NAND4_X1 _21611_ ( .A1(_06595_ ), .A2(_06596_ ), .A3(_06597_ ), .A4(_06602_ ), .ZN(_06603_ ) );
NAND3_X1 _21612_ ( .A1(_06573_ ), .A2(_06592_ ), .A3(_06603_ ), .ZN(_06604_ ) );
BUF_X4 _21613_ ( .A(_06304_ ), .Z(_06605_ ) );
AOI22_X1 _21614_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06605_ ), .B1(_06318_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06606_ ) );
AOI22_X1 _21615_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06321_ ), .B1(_06322_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06607_ ) );
NAND3_X1 _21616_ ( .A1(_06606_ ), .A2(_06320_ ), .A3(_06607_ ), .ZN(_06608_ ) );
BUF_X4 _21617_ ( .A(_06317_ ), .Z(_06609_ ) );
AOI22_X1 _21618_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06605_ ), .B1(_06609_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06610_ ) );
BUF_X4 _21619_ ( .A(_09084_ ), .Z(_06611_ ) );
AOI22_X1 _21620_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06325_ ), .B1(_06327_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06612_ ) );
NAND3_X1 _21621_ ( .A1(_06610_ ), .A2(_06611_ ), .A3(_06612_ ), .ZN(_06613_ ) );
NAND3_X1 _21622_ ( .A1(_06303_ ), .A2(_06608_ ), .A3(_06613_ ), .ZN(_06614_ ) );
NAND3_X1 _21623_ ( .A1(_06604_ ), .A2(_11056_ ), .A3(_06614_ ), .ZN(_06615_ ) );
NAND3_X1 _21624_ ( .A1(_06585_ ), .A2(_10744_ ), .A3(_06615_ ), .ZN(_06616_ ) );
AND3_X1 _21625_ ( .A1(_06456_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06240_ ), .ZN(_06617_ ) );
AOI221_X4 _21626_ ( .A(_06617_ ), .B1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06242_ ), .C1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .C2(_09627_ ), .ZN(_06618_ ) );
BUF_X4 _21627_ ( .A(_09070_ ), .Z(_06619_ ) );
NAND3_X1 _21628_ ( .A1(_06619_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06249_ ), .ZN(_06620_ ) );
NAND3_X1 _21629_ ( .A1(_06618_ ), .A2(_06308_ ), .A3(_06620_ ), .ZN(_06621_ ) );
BUF_X4 _21630_ ( .A(_06326_ ), .Z(_06622_ ) );
AOI22_X1 _21631_ ( .A1(_06342_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06622_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06623_ ) );
OAI211_X1 _21632_ ( .A(_06333_ ), .B(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06600_ ), .C2(_06601_ ), .ZN(_06624_ ) );
BUF_X4 _21633_ ( .A(_06165_ ), .Z(_06625_ ) );
NAND3_X1 _21634_ ( .A1(_06625_ ), .A2(_06331_ ), .A3(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06626_ ) );
NAND3_X1 _21635_ ( .A1(_06623_ ), .A2(_06624_ ), .A3(_06626_ ), .ZN(_06627_ ) );
OAI211_X1 _21636_ ( .A(_06621_ ), .B(_06204_ ), .C1(_06198_ ), .C2(_06627_ ), .ZN(_06628_ ) );
BUF_X4 _21637_ ( .A(_05868_ ), .Z(_06629_ ) );
BUF_X4 _21638_ ( .A(_05869_ ), .Z(_06630_ ) );
OAI211_X1 _21639_ ( .A(_06256_ ), .B(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06629_ ), .C2(_06630_ ), .ZN(_06631_ ) );
INV_X1 _21640_ ( .A(_06631_ ), .ZN(_06632_ ) );
AOI221_X4 _21641_ ( .A(_06632_ ), .B1(_06231_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C2(_09627_ ), .ZN(_06633_ ) );
NAND3_X1 _21642_ ( .A1(_06309_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06590_ ), .ZN(_06634_ ) );
AOI21_X1 _21643_ ( .A(_06192_ ), .B1(_06633_ ), .B2(_06634_ ), .ZN(_06635_ ) );
BUF_X4 _21644_ ( .A(_06157_ ), .Z(_06636_ ) );
BUF_X4 _21645_ ( .A(_09745_ ), .Z(_06637_ ) );
BUF_X4 _21646_ ( .A(_09123_ ), .Z(_06638_ ) );
AOI22_X1 _21647_ ( .A1(_06637_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06638_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06639_ ) );
BUF_X4 _21648_ ( .A(_06212_ ), .Z(_06640_ ) );
AOI22_X1 _21649_ ( .A1(_06343_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06640_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06641_ ) );
AOI21_X1 _21650_ ( .A(_06636_ ), .B1(_06639_ ), .B2(_06641_ ), .ZN(_06642_ ) );
OAI21_X1 _21651_ ( .A(_10050_ ), .B1(_06635_ ), .B2(_06642_ ), .ZN(_06643_ ) );
NAND3_X1 _21652_ ( .A1(_06628_ ), .A2(_10053_ ), .A3(_06643_ ), .ZN(_06644_ ) );
BUF_X4 _21653_ ( .A(_09481_ ), .Z(_06645_ ) );
AOI22_X1 _21654_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06342_ ), .B1(_06263_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06646_ ) );
AOI22_X1 _21655_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06379_ ), .B1(_06380_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06647_ ) );
AOI21_X1 _21656_ ( .A(_06192_ ), .B1(_06646_ ), .B2(_06647_ ), .ZN(_06648_ ) );
BUF_X4 _21657_ ( .A(_06383_ ), .Z(_06649_ ) );
AOI22_X1 _21658_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06421_ ), .B1(_06649_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06650_ ) );
AOI22_X1 _21659_ ( .A1(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06347_ ), .B1(_06640_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06651_ ) );
AOI21_X1 _21660_ ( .A(_06636_ ), .B1(_06650_ ), .B2(_06651_ ), .ZN(_06652_ ) );
OAI21_X1 _21661_ ( .A(_06645_ ), .B1(_06648_ ), .B2(_06652_ ), .ZN(_06653_ ) );
BUF_X4 _21662_ ( .A(_09664_ ), .Z(_06654_ ) );
AOI22_X1 _21663_ ( .A1(_06476_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06470_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06655_ ) );
OAI211_X1 _21664_ ( .A(_06350_ ), .B(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06353_ ), .C2(_06356_ ), .ZN(_06656_ ) );
NAND3_X1 _21665_ ( .A1(_06483_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06484_ ), .ZN(_06657_ ) );
NAND4_X1 _21666_ ( .A1(_06655_ ), .A2(_06192_ ), .A3(_06656_ ), .A4(_06657_ ), .ZN(_06658_ ) );
AOI22_X1 _21667_ ( .A1(_06346_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06220_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06659_ ) );
AOI22_X1 _21668_ ( .A1(_06469_ ), .A2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06380_ ), .B2(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06660_ ) );
NAND3_X1 _21669_ ( .A1(_06659_ ), .A2(_06660_ ), .A3(_06565_ ), .ZN(_06661_ ) );
NAND3_X1 _21670_ ( .A1(_09056_ ), .A2(_06658_ ), .A3(_06661_ ), .ZN(_06662_ ) );
NAND3_X1 _21671_ ( .A1(_06653_ ), .A2(_06654_ ), .A3(_06662_ ), .ZN(_06663_ ) );
NAND3_X1 _21672_ ( .A1(_06644_ ), .A2(_06338_ ), .A3(_06663_ ), .ZN(_06664_ ) );
NAND3_X1 _21673_ ( .A1(_06616_ ), .A2(_09604_ ), .A3(_06664_ ), .ZN(_06665_ ) );
NAND3_X1 _21674_ ( .A1(_06554_ ), .A2(_09035_ ), .A3(_06665_ ), .ZN(_06666_ ) );
AND3_X1 _21675_ ( .A1(_06455_ ), .A2(_06666_ ), .A3(_06077_ ), .ZN(\load_data_out[6] ) );
INV_X1 _21676_ ( .A(\load_data_out[6] ), .ZN(_06667_ ) );
OAI21_X1 _21677_ ( .A(_06667_ ), .B1(_09667_ ), .B2(_06130_ ), .ZN(_06668_ ) );
AOI21_X1 _21678_ ( .A(_06142_ ), .B1(_06668_ ), .B2(_06102_ ), .ZN(_06669_ ) );
NOR2_X1 _21679_ ( .A1(_06669_ ), .A2(_06137_ ), .ZN(_00023_ ) );
OAI22_X1 _21680_ ( .A1(_09888_ ), .A2(_05731_ ), .B1(_09105_ ), .B2(_09061_ ), .ZN(_06670_ ) );
BUF_X4 _21681_ ( .A(_09068_ ), .Z(_06671_ ) );
NAND3_X1 _21682_ ( .A1(_06671_ ), .A2(_09093_ ), .A3(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06672_ ) );
INV_X1 _21683_ ( .A(_06672_ ), .ZN(_06673_ ) );
AOI221_X4 _21684_ ( .A(_06673_ ), .B1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06430_ ), .C1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06212_ ), .ZN(_06674_ ) );
BUF_X4 _21685_ ( .A(_06248_ ), .Z(_06675_ ) );
NAND3_X1 _21686_ ( .A1(_06561_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06675_ ), .ZN(_06676_ ) );
AOI21_X1 _21687_ ( .A(_06596_ ), .B1(_06674_ ), .B2(_06676_ ), .ZN(_06677_ ) );
CLKBUF_X2 _21688_ ( .A(_06018_ ), .Z(_06678_ ) );
NAND3_X1 _21689_ ( .A1(_06145_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06678_ ), .ZN(_06679_ ) );
INV_X1 _21690_ ( .A(_06679_ ), .ZN(_06680_ ) );
AOI221_X4 _21691_ ( .A(_06680_ ), .B1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06178_ ), .C1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06150_ ), .ZN(_06681_ ) );
NAND3_X1 _21692_ ( .A1(_06459_ ), .A2(_06460_ ), .A3(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06682_ ) );
AOI21_X1 _21693_ ( .A(_06514_ ), .B1(_06681_ ), .B2(_06682_ ), .ZN(_06683_ ) );
BUF_X4 _21694_ ( .A(_09055_ ), .Z(_06684_ ) );
NOR3_X1 _21695_ ( .A1(_06677_ ), .A2(_06683_ ), .A3(_06684_ ), .ZN(_06685_ ) );
AND3_X1 _21696_ ( .A1(_06228_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06240_ ), .ZN(_06686_ ) );
AOI221_X4 _21697_ ( .A(_06686_ ), .B1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06242_ ), .C1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06285_ ), .ZN(_06687_ ) );
NAND3_X1 _21698_ ( .A1(_06619_ ), .A2(_06569_ ), .A3(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06688_ ) );
NAND3_X1 _21699_ ( .A1(_06687_ ), .A2(_06556_ ), .A3(_06688_ ), .ZN(_06689_ ) );
AND3_X1 _21700_ ( .A1(_06159_ ), .A2(_06391_ ), .A3(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06690_ ) );
AOI221_X4 _21701_ ( .A(_06690_ ), .B1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06189_ ), .C1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06190_ ), .ZN(_06691_ ) );
NAND3_X1 _21702_ ( .A1(_06246_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06311_ ), .ZN(_06692_ ) );
NAND3_X1 _21703_ ( .A1(_06691_ ), .A2(_06565_ ), .A3(_06692_ ), .ZN(_06693_ ) );
AOI21_X1 _21704_ ( .A(_09482_ ), .B1(_06689_ ), .B2(_06693_ ), .ZN(_06694_ ) );
NOR3_X1 _21705_ ( .A1(_06685_ ), .A2(_06694_ ), .A3(_06654_ ), .ZN(_06695_ ) );
AOI22_X1 _21706_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06605_ ), .B1(_06609_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06696_ ) );
BUF_X4 _21707_ ( .A(_06210_ ), .Z(_06697_ ) );
AOI22_X1 _21708_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06697_ ), .B1(_06360_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06698_ ) );
AOI21_X1 _21709_ ( .A(_06329_ ), .B1(_06696_ ), .B2(_06698_ ), .ZN(_06699_ ) );
BUF_X4 _21710_ ( .A(_06157_ ), .Z(_06700_ ) );
AOI22_X1 _21711_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06637_ ), .B1(_06366_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06701_ ) );
BUF_X4 _21712_ ( .A(_06212_ ), .Z(_06702_ ) );
AOI22_X1 _21713_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06369_ ), .B1(_06702_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06703_ ) );
AOI21_X1 _21714_ ( .A(_06700_ ), .B1(_06701_ ), .B2(_06703_ ), .ZN(_06704_ ) );
OAI21_X1 _21715_ ( .A(_06315_ ), .B1(_06699_ ), .B2(_06704_ ), .ZN(_06705_ ) );
AOI22_X1 _21716_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06605_ ), .B1(_06318_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06706_ ) );
AOI22_X1 _21717_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06321_ ), .B1(_06360_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06707_ ) );
NAND3_X1 _21718_ ( .A1(_06706_ ), .A2(_06320_ ), .A3(_06707_ ), .ZN(_06708_ ) );
AOI22_X1 _21719_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06346_ ), .B1(_06609_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06709_ ) );
AOI22_X1 _21720_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06325_ ), .B1(_06327_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06710_ ) );
NAND3_X1 _21721_ ( .A1(_06709_ ), .A2(_06611_ ), .A3(_06710_ ), .ZN(_06711_ ) );
NAND3_X1 _21722_ ( .A1(_06303_ ), .A2(_06708_ ), .A3(_06711_ ), .ZN(_06712_ ) );
AOI21_X1 _21723_ ( .A(_09594_ ), .B1(_06705_ ), .B2(_06712_ ), .ZN(_06713_ ) );
OAI21_X1 _21724_ ( .A(_09489_ ), .B1(_06695_ ), .B2(_06713_ ), .ZN(_06714_ ) );
AND3_X1 _21725_ ( .A1(_06439_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06146_ ), .ZN(_06715_ ) );
BUF_X4 _21726_ ( .A(_09528_ ), .Z(_06716_ ) );
AOI221_X4 _21727_ ( .A(_06715_ ), .B1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06716_ ), .C1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06298_ ), .ZN(_06717_ ) );
BUF_X4 _21728_ ( .A(_09070_ ), .Z(_06718_ ) );
NAND3_X1 _21729_ ( .A1(_06718_ ), .A2(_09095_ ), .A3(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06719_ ) );
NAND3_X1 _21730_ ( .A1(_06717_ ), .A2(_06576_ ), .A3(_06719_ ), .ZN(_06720_ ) );
BUF_X4 _21731_ ( .A(_06255_ ), .Z(_06721_ ) );
BUF_X4 _21732_ ( .A(_06229_ ), .Z(_06722_ ) );
MUX2_X1 _21733_ ( .A(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .S(_06722_ ), .Z(_06723_ ) );
MUX2_X1 _21734_ ( .A(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .S(_06543_ ), .Z(_06724_ ) );
BUF_X4 _21735_ ( .A(_06440_ ), .Z(_06725_ ) );
MUX2_X1 _21736_ ( .A(_06723_ ), .B(_06724_ ), .S(_06725_ ), .Z(_06726_ ) );
OAI211_X1 _21737_ ( .A(_06720_ ), .B(_06303_ ), .C1(_06721_ ), .C2(_06726_ ), .ZN(_06727_ ) );
NAND3_X1 _21738_ ( .A1(_06671_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06399_ ), .ZN(_06728_ ) );
INV_X1 _21739_ ( .A(_06728_ ), .ZN(_06729_ ) );
AOI221_X4 _21740_ ( .A(_06729_ ), .B1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06430_ ), .C1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06326_ ), .ZN(_06730_ ) );
NAND3_X1 _21741_ ( .A1(_06561_ ), .A2(_06562_ ), .A3(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06731_ ) );
AOI21_X1 _21742_ ( .A(_06245_ ), .B1(_06730_ ), .B2(_06731_ ), .ZN(_06732_ ) );
OAI211_X1 _21743_ ( .A(_06229_ ), .B(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06629_ ), .C2(_06630_ ), .ZN(_06733_ ) );
INV_X1 _21744_ ( .A(_06733_ ), .ZN(_06734_ ) );
AOI221_X4 _21745_ ( .A(_06734_ ), .B1(_06716_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C2(_06383_ ), .ZN(_06735_ ) );
BUF_X4 _21746_ ( .A(_06248_ ), .Z(_06736_ ) );
NAND3_X1 _21747_ ( .A1(_06619_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06736_ ), .ZN(_06737_ ) );
AOI21_X1 _21748_ ( .A(_06219_ ), .B1(_06735_ ), .B2(_06737_ ), .ZN(_06738_ ) );
OAI21_X1 _21749_ ( .A(_10261_ ), .B1(_06732_ ), .B2(_06738_ ), .ZN(_06739_ ) );
NAND3_X1 _21750_ ( .A1(_06727_ ), .A2(_11056_ ), .A3(_06739_ ), .ZN(_06740_ ) );
BUF_X4 _21751_ ( .A(_06504_ ), .Z(_06741_ ) );
AOI22_X1 _21752_ ( .A1(_06741_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06321_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06742_ ) );
BUF_X4 _21753_ ( .A(_06352_ ), .Z(_06743_ ) );
BUF_X4 _21754_ ( .A(_06355_ ), .Z(_06744_ ) );
OAI211_X1 _21755_ ( .A(_06460_ ), .B(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06743_ ), .C2(_06744_ ), .ZN(_06745_ ) );
NAND3_X1 _21756_ ( .A1(_06568_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06736_ ), .ZN(_06746_ ) );
NAND4_X1 _21757_ ( .A1(_06742_ ), .A2(_06234_ ), .A3(_06745_ ), .A4(_06746_ ), .ZN(_06747_ ) );
AOI22_X1 _21758_ ( .A1(_06580_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06697_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06748_ ) );
OAI211_X1 _21759_ ( .A(_06331_ ), .B(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06587_ ), .C2(_06588_ ), .ZN(_06749_ ) );
NAND3_X1 _21760_ ( .A1(_06619_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06249_ ), .ZN(_06750_ ) );
NAND4_X1 _21761_ ( .A1(_06748_ ), .A2(_06320_ ), .A3(_06749_ ), .A4(_06750_ ), .ZN(_06751_ ) );
NAND3_X1 _21762_ ( .A1(_10261_ ), .A2(_06747_ ), .A3(_06751_ ), .ZN(_06752_ ) );
AOI22_X1 _21763_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06305_ ), .B1(_06469_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06753_ ) );
AOI22_X1 _21764_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06339_ ), .B1(_06340_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06754_ ) );
NAND3_X1 _21765_ ( .A1(_06753_ ), .A2(_06582_ ), .A3(_06754_ ), .ZN(_06755_ ) );
AOI22_X1 _21766_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06305_ ), .B1(_06469_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06756_ ) );
BUF_X4 _21767_ ( .A(_06179_ ), .Z(_06757_ ) );
AOI22_X1 _21768_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06757_ ), .B1(_06306_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06758_ ) );
NAND3_X1 _21769_ ( .A1(_06756_ ), .A2(_06576_ ), .A3(_06758_ ), .ZN(_06759_ ) );
NAND3_X1 _21770_ ( .A1(_06555_ ), .A2(_06755_ ), .A3(_06759_ ), .ZN(_06760_ ) );
NAND3_X1 _21771_ ( .A1(_06752_ ), .A2(_09784_ ), .A3(_06760_ ), .ZN(_06761_ ) );
NAND3_X1 _21772_ ( .A1(_06740_ ), .A2(_06143_ ), .A3(_06761_ ), .ZN(_06762_ ) );
NAND3_X1 _21773_ ( .A1(_06714_ ), .A2(_09491_ ), .A3(_06762_ ), .ZN(_06763_ ) );
AND3_X1 _21774_ ( .A1(_06439_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06296_ ), .ZN(_06764_ ) );
AOI221_X4 _21775_ ( .A(_06764_ ), .B1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06163_ ), .C1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06298_ ), .ZN(_06765_ ) );
NAND3_X1 _21776_ ( .A1(_06718_ ), .A2(_09095_ ), .A3(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06766_ ) );
NAND3_X1 _21777_ ( .A1(_06765_ ), .A2(_06300_ ), .A3(_06766_ ), .ZN(_06767_ ) );
AOI22_X1 _21778_ ( .A1(_06316_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06306_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06768_ ) );
NAND3_X1 _21779_ ( .A1(_06152_ ), .A2(_06154_ ), .A3(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06769_ ) );
NAND3_X1 _21780_ ( .A1(_06246_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06311_ ), .ZN(_06770_ ) );
NAND4_X1 _21781_ ( .A1(_06768_ ), .A2(_06308_ ), .A3(_06769_ ), .A4(_06770_ ), .ZN(_06771_ ) );
NAND3_X1 _21782_ ( .A1(_06767_ ), .A2(_06303_ ), .A3(_06771_ ), .ZN(_06772_ ) );
AOI22_X1 _21783_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06316_ ), .B1(_06318_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06773_ ) );
AOI22_X1 _21784_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06757_ ), .B1(_06322_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06774_ ) );
NAND3_X1 _21785_ ( .A1(_06773_ ), .A2(_06234_ ), .A3(_06774_ ), .ZN(_06775_ ) );
AOI22_X1 _21786_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06757_ ), .B1(_06340_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06776_ ) );
AOI22_X1 _21787_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06365_ ), .B1(_06263_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06777_ ) );
NAND3_X1 _21788_ ( .A1(_06776_ ), .A2(_06245_ ), .A3(_06777_ ), .ZN(_06778_ ) );
NAND3_X1 _21789_ ( .A1(_06315_ ), .A2(_06775_ ), .A3(_06778_ ), .ZN(_06779_ ) );
AOI21_X1 _21790_ ( .A(_09487_ ), .B1(_06772_ ), .B2(_06779_ ), .ZN(_06780_ ) );
BUF_X4 _21791_ ( .A(_06317_ ), .Z(_06781_ ) );
AOI22_X1 _21792_ ( .A1(_06781_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06347_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06782_ ) );
BUF_X4 _21793_ ( .A(_06248_ ), .Z(_06783_ ) );
NAND3_X1 _21794_ ( .A1(_06330_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06783_ ), .ZN(_06784_ ) );
OAI211_X1 _21795_ ( .A(_06350_ ), .B(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06353_ ), .C2(_06356_ ), .ZN(_06785_ ) );
NAND4_X1 _21796_ ( .A1(_06782_ ), .A2(_06209_ ), .A3(_06784_ ), .A4(_06785_ ), .ZN(_06786_ ) );
AOI22_X1 _21797_ ( .A1(_06316_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06594_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06787_ ) );
AOI22_X1 _21798_ ( .A1(_06781_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06327_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06788_ ) );
NAND3_X1 _21799_ ( .A1(_06787_ ), .A2(_06788_ ), .A3(_06362_ ), .ZN(_06789_ ) );
NAND3_X1 _21800_ ( .A1(_06315_ ), .A2(_06786_ ), .A3(_06789_ ), .ZN(_06790_ ) );
AOI22_X1 _21801_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06342_ ), .B1(_06263_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06791_ ) );
AOI22_X1 _21802_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06594_ ), .B1(_06370_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06792_ ) );
NAND3_X1 _21803_ ( .A1(_06791_ ), .A2(_06368_ ), .A3(_06792_ ), .ZN(_06793_ ) );
BUF_X4 _21804_ ( .A(_06210_ ), .Z(_06794_ ) );
AOI22_X1 _21805_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06794_ ), .B1(_06274_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06795_ ) );
NAND3_X1 _21806_ ( .A1(_06483_ ), .A2(_06167_ ), .A3(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06796_ ) );
BUF_X4 _21807_ ( .A(_06399_ ), .Z(_06797_ ) );
BUF_X4 _21808_ ( .A(_06797_ ), .Z(_06798_ ) );
NAND3_X1 _21809_ ( .A1(_06166_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06798_ ), .ZN(_06799_ ) );
NAND4_X1 _21810_ ( .A1(_06795_ ), .A2(_06514_ ), .A3(_06796_ ), .A4(_06799_ ), .ZN(_06800_ ) );
NAND3_X1 _21811_ ( .A1(_09056_ ), .A2(_06793_ ), .A3(_06800_ ), .ZN(_06801_ ) );
AOI21_X1 _21812_ ( .A(_09665_ ), .B1(_06790_ ), .B2(_06801_ ), .ZN(_06802_ ) );
OAI21_X1 _21813_ ( .A(_06143_ ), .B1(_06780_ ), .B2(_06802_ ), .ZN(_06803_ ) );
NAND3_X1 _21814_ ( .A1(_06671_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06399_ ), .ZN(_06804_ ) );
INV_X1 _21815_ ( .A(_06804_ ), .ZN(_06805_ ) );
AOI221_X4 _21816_ ( .A(_06805_ ), .B1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06259_ ), .C1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C2(_06317_ ), .ZN(_06806_ ) );
NAND3_X1 _21817_ ( .A1(_10432_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06675_ ), .ZN(_06807_ ) );
NAND3_X1 _21818_ ( .A1(_06806_ ), .A2(_06300_ ), .A3(_06807_ ), .ZN(_06808_ ) );
AOI22_X1 _21819_ ( .A1(_06574_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_09530_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06809_ ) );
NAND3_X1 _21820_ ( .A1(_06246_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06736_ ), .ZN(_06810_ ) );
BUF_X4 _21821_ ( .A(_06153_ ), .Z(_06811_ ) );
NAND3_X1 _21822_ ( .A1(_06619_ ), .A2(_06811_ ), .A3(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06812_ ) );
NAND4_X1 _21823_ ( .A1(_06809_ ), .A2(_06234_ ), .A3(_06810_ ), .A4(_06812_ ), .ZN(_06813_ ) );
NAND3_X1 _21824_ ( .A1(_06808_ ), .A2(_06555_ ), .A3(_06813_ ), .ZN(_06814_ ) );
AOI22_X1 _21825_ ( .A1(_06580_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06594_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06815_ ) );
NAND3_X1 _21826_ ( .A1(_06309_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06590_ ), .ZN(_06816_ ) );
OAI211_X1 _21827_ ( .A(_06599_ ), .B(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06587_ ), .C2(_06588_ ), .ZN(_06817_ ) );
NAND4_X1 _21828_ ( .A1(_06815_ ), .A2(_06308_ ), .A3(_06816_ ), .A4(_06817_ ), .ZN(_06818_ ) );
AOI22_X1 _21829_ ( .A1(_06574_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06697_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06819_ ) );
AOI22_X1 _21830_ ( .A1(_06580_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06306_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06820_ ) );
NAND3_X1 _21831_ ( .A1(_06819_ ), .A2(_06820_ ), .A3(_06320_ ), .ZN(_06821_ ) );
NAND3_X1 _21832_ ( .A1(_06573_ ), .A2(_06818_ ), .A3(_06821_ ), .ZN(_06822_ ) );
NAND3_X1 _21833_ ( .A1(_06814_ ), .A2(_10053_ ), .A3(_06822_ ), .ZN(_06823_ ) );
AOI22_X1 _21834_ ( .A1(_06593_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06594_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06824_ ) );
OAI211_X1 _21835_ ( .A(_06515_ ), .B(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06587_ ), .C2(_06588_ ), .ZN(_06825_ ) );
NAND3_X1 _21836_ ( .A1(_06459_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06311_ ), .ZN(_06826_ ) );
NAND4_X1 _21837_ ( .A1(_06824_ ), .A2(_06308_ ), .A3(_06825_ ), .A4(_06826_ ), .ZN(_06827_ ) );
AOI22_X1 _21838_ ( .A1(_06593_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06369_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06828_ ) );
NAND3_X1 _21839_ ( .A1(_06459_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06590_ ), .ZN(_06829_ ) );
OAI211_X1 _21840_ ( .A(_06599_ ), .B(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06600_ ), .C2(_06601_ ), .ZN(_06830_ ) );
NAND4_X1 _21841_ ( .A1(_06828_ ), .A2(_06596_ ), .A3(_06829_ ), .A4(_06830_ ), .ZN(_06831_ ) );
NAND3_X1 _21842_ ( .A1(_06573_ ), .A2(_06827_ ), .A3(_06831_ ), .ZN(_06832_ ) );
AOI22_X1 _21843_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06757_ ), .B1(_06306_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06833_ ) );
AOI22_X1 _21844_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06365_ ), .B1(_06263_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06834_ ) );
NAND3_X1 _21845_ ( .A1(_06833_ ), .A2(_06611_ ), .A3(_06834_ ), .ZN(_06835_ ) );
BUF_X4 _21846_ ( .A(_06317_ ), .Z(_06836_ ) );
AOI22_X1 _21847_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06346_ ), .B1(_06836_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06837_ ) );
AOI22_X1 _21848_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06325_ ), .B1(_06622_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06838_ ) );
NAND3_X1 _21849_ ( .A1(_06837_ ), .A2(_06245_ ), .A3(_06838_ ), .ZN(_06839_ ) );
NAND3_X1 _21850_ ( .A1(_06303_ ), .A2(_06835_ ), .A3(_06839_ ), .ZN(_06840_ ) );
NAND3_X1 _21851_ ( .A1(_06832_ ), .A2(_11056_ ), .A3(_06840_ ), .ZN(_06841_ ) );
NAND3_X1 _21852_ ( .A1(_06823_ ), .A2(_10744_ ), .A3(_06841_ ), .ZN(_06842_ ) );
NAND3_X1 _21853_ ( .A1(_06803_ ), .A2(_02457_ ), .A3(_06842_ ), .ZN(_06843_ ) );
NAND3_X1 _21854_ ( .A1(_06763_ ), .A2(_09493_ ), .A3(_06843_ ), .ZN(_06844_ ) );
AND3_X1 _21855_ ( .A1(_06557_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06678_ ), .ZN(_06845_ ) );
AOI221_X4 _21856_ ( .A(_06845_ ), .B1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06559_ ), .C1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06232_ ), .ZN(_06846_ ) );
NAND3_X1 _21857_ ( .A1(_06235_ ), .A2(_06236_ ), .A3(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06847_ ) );
NAND3_X1 _21858_ ( .A1(_06846_ ), .A2(_06234_ ), .A3(_06847_ ), .ZN(_06848_ ) );
AND3_X1 _21859_ ( .A1(_06239_ ), .A2(_06391_ ), .A3(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06849_ ) );
AOI221_X4 _21860_ ( .A(_06849_ ), .B1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06242_ ), .C1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06285_ ), .ZN(_06850_ ) );
NAND3_X1 _21861_ ( .A1(_06246_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06249_ ), .ZN(_06851_ ) );
NAND3_X1 _21862_ ( .A1(_06850_ ), .A2(_06245_ ), .A3(_06851_ ), .ZN(_06852_ ) );
NAND3_X1 _21863_ ( .A1(_06848_ ), .A2(_06852_ ), .A3(_06252_ ), .ZN(_06853_ ) );
AOI22_X1 _21864_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06365_ ), .B1(_06366_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06854_ ) );
AOI22_X1 _21865_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06369_ ), .B1(_06370_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06855_ ) );
NAND3_X1 _21866_ ( .A1(_06854_ ), .A2(_06368_ ), .A3(_06855_ ), .ZN(_06856_ ) );
BUF_X4 _21867_ ( .A(_09745_ ), .Z(_06857_ ) );
AOI22_X1 _21868_ ( .A1(_06857_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06347_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06858_ ) );
AOI22_X1 _21869_ ( .A1(_06476_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06370_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06859_ ) );
NAND3_X1 _21870_ ( .A1(_06858_ ), .A2(_06859_ ), .A3(_06219_ ), .ZN(_06860_ ) );
NAND3_X1 _21871_ ( .A1(_06645_ ), .A2(_06856_ ), .A3(_06860_ ), .ZN(_06861_ ) );
AOI21_X1 _21872_ ( .A(_09665_ ), .B1(_06853_ ), .B2(_06861_ ), .ZN(_06862_ ) );
AOI22_X1 _21873_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_09746_ ), .B1(_06540_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06863_ ) );
BUF_X4 _21874_ ( .A(_06424_ ), .Z(_06864_ ) );
AOI22_X1 _21875_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06470_ ), .B1(_06864_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06865_ ) );
AOI21_X1 _21876_ ( .A(_06405_ ), .B1(_06863_ ), .B2(_06865_ ), .ZN(_06866_ ) );
AOI22_X1 _21877_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06444_ ), .B1(_06527_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06867_ ) );
AOI22_X1 _21878_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06422_ ), .B1(_06268_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06868_ ) );
AOI21_X1 _21879_ ( .A(_06433_ ), .B1(_06867_ ), .B2(_06868_ ), .ZN(_06869_ ) );
OAI21_X1 _21880_ ( .A(_06463_ ), .B1(_06866_ ), .B2(_06869_ ), .ZN(_06870_ ) );
AOI22_X1 _21881_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06421_ ), .B1(_06429_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06871_ ) );
BUF_X4 _21882_ ( .A(_09123_ ), .Z(_06872_ ) );
AOI22_X1 _21883_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06872_ ), .B1(_06864_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06873_ ) );
NAND3_X1 _21884_ ( .A1(_06871_ ), .A2(_06479_ ), .A3(_06873_ ), .ZN(_06874_ ) );
AOI22_X1 _21885_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06382_ ), .B1(_06540_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06875_ ) );
AOI22_X1 _21886_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06470_ ), .B1(_06425_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06876_ ) );
NAND3_X1 _21887_ ( .A1(_06875_ ), .A2(_06514_ ), .A3(_06876_ ), .ZN(_06877_ ) );
NAND3_X1 _21888_ ( .A1(_06388_ ), .A2(_06874_ ), .A3(_06877_ ), .ZN(_06878_ ) );
AOI21_X1 _21889_ ( .A(_06186_ ), .B1(_06870_ ), .B2(_06878_ ), .ZN(_06879_ ) );
OAI21_X1 _21890_ ( .A(_06227_ ), .B1(_06862_ ), .B2(_06879_ ), .ZN(_06880_ ) );
AND3_X1 _21891_ ( .A1(_06439_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06296_ ), .ZN(_06881_ ) );
AOI221_X4 _21892_ ( .A(_06881_ ), .B1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06716_ ), .C1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06298_ ), .ZN(_06882_ ) );
NAND3_X1 _21893_ ( .A1(_06718_ ), .A2(_09095_ ), .A3(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06883_ ) );
NAND3_X1 _21894_ ( .A1(_06882_ ), .A2(_06576_ ), .A3(_06883_ ), .ZN(_06884_ ) );
AND3_X1 _21895_ ( .A1(_06557_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06678_ ), .ZN(_06885_ ) );
AOI221_X4 _21896_ ( .A(_06885_ ), .B1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06559_ ), .C1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06232_ ), .ZN(_06886_ ) );
NAND3_X1 _21897_ ( .A1(_06235_ ), .A2(_06236_ ), .A3(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06887_ ) );
NAND3_X1 _21898_ ( .A1(_06886_ ), .A2(_06582_ ), .A3(_06887_ ), .ZN(_06888_ ) );
NAND3_X1 _21899_ ( .A1(_06884_ ), .A2(_06888_ ), .A3(_10050_ ), .ZN(_06889_ ) );
BUF_X4 _21900_ ( .A(_09481_ ), .Z(_06890_ ) );
AOI22_X1 _21901_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06346_ ), .B1(_06836_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06891_ ) );
AOI22_X1 _21902_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06325_ ), .B1(_06622_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06892_ ) );
NAND3_X1 _21903_ ( .A1(_06891_ ), .A2(_06556_ ), .A3(_06892_ ), .ZN(_06893_ ) );
AOI22_X1 _21904_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06857_ ), .B1(_06343_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06894_ ) );
AOI22_X1 _21905_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06379_ ), .B1(_06622_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06895_ ) );
NAND3_X1 _21906_ ( .A1(_06894_ ), .A2(_06596_ ), .A3(_06895_ ), .ZN(_06896_ ) );
NAND3_X1 _21907_ ( .A1(_06890_ ), .A2(_06893_ ), .A3(_06896_ ), .ZN(_06897_ ) );
NAND3_X1 _21908_ ( .A1(_06889_ ), .A2(_09487_ ), .A3(_06897_ ), .ZN(_06898_ ) );
NAND3_X1 _21909_ ( .A1(_06145_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06146_ ), .ZN(_06899_ ) );
INV_X1 _21910_ ( .A(_06899_ ), .ZN(_06900_ ) );
AOI221_X4 _21911_ ( .A(_06900_ ), .B1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06149_ ), .C1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06150_ ), .ZN(_06901_ ) );
NAND3_X1 _21912_ ( .A1(_06152_ ), .A2(_06154_ ), .A3(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06902_ ) );
AOI21_X1 _21913_ ( .A(_06144_ ), .B1(_06901_ ), .B2(_06902_ ), .ZN(_06903_ ) );
NAND3_X1 _21914_ ( .A1(_06239_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06256_ ), .ZN(_06904_ ) );
INV_X1 _21915_ ( .A(_06904_ ), .ZN(_06905_ ) );
AOI221_X4 _21916_ ( .A(_06905_ ), .B1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06178_ ), .C1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06259_ ), .ZN(_06906_ ) );
NAND3_X1 _21917_ ( .A1(_06193_ ), .A2(_06194_ ), .A3(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06907_ ) );
AOI21_X1 _21918_ ( .A(_06636_ ), .B1(_06906_ ), .B2(_06907_ ), .ZN(_06908_ ) );
OAI21_X1 _21919_ ( .A(_06645_ ), .B1(_06903_ ), .B2(_06908_ ), .ZN(_06909_ ) );
AOI22_X1 _21920_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06421_ ), .B1(_06649_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06910_ ) );
AOI22_X1 _21921_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06347_ ), .B1(_06640_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06911_ ) );
AOI21_X1 _21922_ ( .A(_06255_ ), .B1(_06910_ ), .B2(_06911_ ), .ZN(_06912_ ) );
AOI22_X1 _21923_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06267_ ), .B1(_09795_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06913_ ) );
BUF_X4 _21924_ ( .A(_09123_ ), .Z(_06914_ ) );
BUF_X4 _21925_ ( .A(_06150_ ), .Z(_06915_ ) );
AOI22_X1 _21926_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06914_ ), .B1(_06915_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06916_ ) );
AOI21_X1 _21927_ ( .A(_06158_ ), .B1(_06913_ ), .B2(_06916_ ), .ZN(_06917_ ) );
OAI21_X1 _21928_ ( .A(_06684_ ), .B1(_06912_ ), .B2(_06917_ ), .ZN(_06918_ ) );
NAND3_X1 _21929_ ( .A1(_06909_ ), .A2(_06654_ ), .A3(_06918_ ), .ZN(_06919_ ) );
NAND3_X1 _21930_ ( .A1(_06898_ ), .A2(_06919_ ), .A3(_06338_ ), .ZN(_06920_ ) );
AOI21_X1 _21931_ ( .A(_02457_ ), .B1(_06880_ ), .B2(_06920_ ), .ZN(_06921_ ) );
AND3_X1 _21932_ ( .A1(_06456_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06240_ ), .ZN(_06922_ ) );
BUF_X4 _21933_ ( .A(_05865_ ), .Z(_06923_ ) );
AOI221_X4 _21934_ ( .A(_06922_ ), .B1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06923_ ), .C1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06176_ ), .ZN(_06924_ ) );
BUF_X4 _21935_ ( .A(_09070_ ), .Z(_06925_ ) );
NAND3_X1 _21936_ ( .A1(_06925_ ), .A2(_06811_ ), .A3(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06926_ ) );
NAND3_X1 _21937_ ( .A1(_06924_ ), .A2(_06596_ ), .A3(_06926_ ), .ZN(_06927_ ) );
AOI22_X1 _21938_ ( .A1(_06421_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06221_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06928_ ) );
BUF_X4 _21939_ ( .A(_09119_ ), .Z(_06929_ ) );
NAND3_X1 _21940_ ( .A1(_06166_ ), .A2(_06167_ ), .A3(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06930_ ) );
BUF_X4 _21941_ ( .A(_06797_ ), .Z(_06931_ ) );
NAND3_X1 _21942_ ( .A1(_06725_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06931_ ), .ZN(_06932_ ) );
NAND4_X1 _21943_ ( .A1(_06928_ ), .A2(_06929_ ), .A3(_06930_ ), .A4(_06932_ ), .ZN(_06933_ ) );
NAND3_X1 _21944_ ( .A1(_06927_ ), .A2(_06684_ ), .A3(_06933_ ), .ZN(_06934_ ) );
AOI22_X1 _21945_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_09746_ ), .B1(_06429_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06935_ ) );
AOI22_X1 _21946_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06872_ ), .B1(_06864_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06936_ ) );
NAND3_X1 _21947_ ( .A1(_06935_ ), .A2(_06144_ ), .A3(_06936_ ), .ZN(_06937_ ) );
AOI22_X1 _21948_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06477_ ), .B1(_06425_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06938_ ) );
BUF_X4 _21949_ ( .A(_06598_ ), .Z(_06939_ ) );
NAND3_X1 _21950_ ( .A1(_06398_ ), .A2(_06939_ ), .A3(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06940_ ) );
NAND3_X1 _21951_ ( .A1(_06407_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06408_ ), .ZN(_06941_ ) );
NAND4_X1 _21952_ ( .A1(_06938_ ), .A2(_06390_ ), .A3(_06940_ ), .A4(_06941_ ), .ZN(_06942_ ) );
NAND3_X1 _21953_ ( .A1(_06463_ ), .A2(_06937_ ), .A3(_06942_ ), .ZN(_06943_ ) );
AOI21_X1 _21954_ ( .A(_06186_ ), .B1(_06934_ ), .B2(_06943_ ), .ZN(_06944_ ) );
AOI22_X1 _21955_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06220_ ), .B1(_06213_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06945_ ) );
AOI22_X1 _21956_ ( .A1(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06444_ ), .B1(_06527_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06946_ ) );
NAND3_X1 _21957_ ( .A1(_06945_ ), .A2(_06514_ ), .A3(_06946_ ), .ZN(_06947_ ) );
AOI22_X1 _21958_ ( .A1(_06421_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_09484_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06948_ ) );
AOI22_X1 _21959_ ( .A1(_06366_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06425_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06949_ ) );
BUF_X4 _21960_ ( .A(_06157_ ), .Z(_06950_ ) );
NAND3_X1 _21961_ ( .A1(_06948_ ), .A2(_06949_ ), .A3(_06950_ ), .ZN(_06951_ ) );
NAND3_X1 _21962_ ( .A1(_06463_ ), .A2(_06947_ ), .A3(_06951_ ), .ZN(_06952_ ) );
AOI22_X1 _21963_ ( .A1(_06429_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06445_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06953_ ) );
NAND3_X1 _21964_ ( .A1(_06407_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06437_ ), .ZN(_06954_ ) );
OAI211_X1 _21965_ ( .A(_06544_ ), .B(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06417_ ), .C2(_06418_ ), .ZN(_06955_ ) );
NAND4_X1 _21966_ ( .A1(_06953_ ), .A2(_06158_ ), .A3(_06954_ ), .A4(_06955_ ), .ZN(_06956_ ) );
AOI22_X1 _21967_ ( .A1(_06522_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06264_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06957_ ) );
AOI22_X1 _21968_ ( .A1(_06649_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06268_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06958_ ) );
NAND3_X1 _21969_ ( .A1(_06957_ ), .A2(_06958_ ), .A3(_06405_ ), .ZN(_06959_ ) );
NAND3_X1 _21970_ ( .A1(_09463_ ), .A2(_06956_ ), .A3(_06959_ ), .ZN(_06960_ ) );
AOI21_X1 _21971_ ( .A(_06413_ ), .B1(_06952_ ), .B2(_06960_ ), .ZN(_06961_ ) );
OAI21_X1 _21972_ ( .A(_06338_ ), .B1(_06944_ ), .B2(_06961_ ), .ZN(_06962_ ) );
AOI22_X1 _21973_ ( .A1(_06469_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06872_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06963_ ) );
BUF_X4 _21974_ ( .A(_09483_ ), .Z(_06964_ ) );
OAI211_X1 _21975_ ( .A(_06350_ ), .B(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06353_ ), .C2(_06356_ ), .ZN(_06965_ ) );
NAND3_X1 _21976_ ( .A1(_06473_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06333_ ), .ZN(_06966_ ) );
NAND4_X1 _21977_ ( .A1(_06963_ ), .A2(_06964_ ), .A3(_06965_ ), .A4(_06966_ ), .ZN(_06967_ ) );
AOI22_X1 _21978_ ( .A1(_06593_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06794_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06968_ ) );
AOI22_X1 _21979_ ( .A1(_06857_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06622_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06969_ ) );
NAND3_X1 _21980_ ( .A1(_06968_ ), .A2(_06969_ ), .A3(_06368_ ), .ZN(_06970_ ) );
NAND3_X1 _21981_ ( .A1(_06890_ ), .A2(_06967_ ), .A3(_06970_ ), .ZN(_06971_ ) );
AOI22_X1 _21982_ ( .A1(_06609_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06914_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06972_ ) );
BUF_X4 _21983_ ( .A(_06157_ ), .Z(_06973_ ) );
OAI211_X1 _21984_ ( .A(_06939_ ), .B(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06480_ ), .C2(_06481_ ), .ZN(_06974_ ) );
NAND3_X1 _21985_ ( .A1(_06492_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06931_ ), .ZN(_06975_ ) );
NAND4_X1 _21986_ ( .A1(_06972_ ), .A2(_06973_ ), .A3(_06974_ ), .A4(_06975_ ), .ZN(_06976_ ) );
AOI22_X1 _21987_ ( .A1(_06836_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_09484_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06977_ ) );
BUF_X4 _21988_ ( .A(_06598_ ), .Z(_06978_ ) );
OAI211_X1 _21989_ ( .A(_06978_ ), .B(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06394_ ), .C2(_06395_ ), .ZN(_06979_ ) );
NAND3_X1 _21990_ ( .A1(_06492_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06931_ ), .ZN(_06980_ ) );
NAND4_X1 _21991_ ( .A1(_06977_ ), .A2(_06929_ ), .A3(_06979_ ), .A4(_06980_ ), .ZN(_06981_ ) );
NAND3_X1 _21992_ ( .A1(_06252_ ), .A2(_06976_ ), .A3(_06981_ ), .ZN(_06982_ ) );
NAND3_X1 _21993_ ( .A1(_06971_ ), .A2(_11196_ ), .A3(_06982_ ), .ZN(_06983_ ) );
AOI22_X1 _21994_ ( .A1(_06318_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06638_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06984_ ) );
NAND3_X1 _21995_ ( .A1(_06166_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06484_ ), .ZN(_06985_ ) );
OAI211_X1 _21996_ ( .A(_06939_ ), .B(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06480_ ), .C2(_06481_ ), .ZN(_06986_ ) );
NAND4_X1 _21997_ ( .A1(_06984_ ), .A2(_06700_ ), .A3(_06985_ ), .A4(_06986_ ), .ZN(_06987_ ) );
AOI22_X1 _21998_ ( .A1(_06857_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06872_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06988_ ) );
AOI22_X1 _21999_ ( .A1(_06476_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06702_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06989_ ) );
NAND3_X1 _22000_ ( .A1(_06988_ ), .A2(_06989_ ), .A3(_06219_ ), .ZN(_06990_ ) );
NAND3_X1 _22001_ ( .A1(_06204_ ), .A2(_06987_ ), .A3(_06990_ ), .ZN(_06991_ ) );
AOI22_X1 _22002_ ( .A1(_06263_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06264_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_06992_ ) );
NAND3_X1 _22003_ ( .A1(_06398_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06931_ ), .ZN(_06993_ ) );
NAND3_X1 _22004_ ( .A1(_06725_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06939_ ), .ZN(_06994_ ) );
NAND4_X1 _22005_ ( .A1(_06992_ ), .A2(_06636_ ), .A3(_06993_ ), .A4(_06994_ ), .ZN(_06995_ ) );
AOI22_X1 _22006_ ( .A1(_06382_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06425_ ), .B2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06996_ ) );
NAND3_X1 _22007_ ( .A1(_06398_ ), .A2(_06350_ ), .A3(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_06997_ ) );
NAND3_X1 _22008_ ( .A1(_06725_ ), .A2(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06401_ ), .ZN(_06998_ ) );
NAND4_X1 _22009_ ( .A1(_06996_ ), .A2(_06405_ ), .A3(_06997_ ), .A4(_06998_ ), .ZN(_06999_ ) );
NAND3_X1 _22010_ ( .A1(_06684_ ), .A2(_06995_ ), .A3(_06999_ ), .ZN(_07000_ ) );
NAND3_X1 _22011_ ( .A1(_06991_ ), .A2(_09594_ ), .A3(_07000_ ), .ZN(_07001_ ) );
NAND3_X1 _22012_ ( .A1(_06983_ ), .A2(_07001_ ), .A3(_06227_ ), .ZN(_07002_ ) );
AOI21_X1 _22013_ ( .A(_09604_ ), .B1(_06962_ ), .B2(_07002_ ), .ZN(_07003_ ) );
OAI21_X1 _22014_ ( .A(_09035_ ), .B1(_06921_ ), .B2(_07003_ ), .ZN(_07004_ ) );
AND3_X1 _22015_ ( .A1(_06844_ ), .A2(_07004_ ), .A3(_06077_ ), .ZN(\load_data_out[5] ) );
INV_X1 _22016_ ( .A(\load_data_out[5] ), .ZN(_07005_ ) );
OAI21_X1 _22017_ ( .A(_07005_ ), .B1(_09888_ ), .B2(_06130_ ), .ZN(_07006_ ) );
AOI21_X1 _22018_ ( .A(_06670_ ), .B1(_07006_ ), .B2(_06102_ ), .ZN(_07007_ ) );
NOR2_X1 _22019_ ( .A1(_07007_ ), .A2(_06137_ ), .ZN(_00024_ ) );
BUF_X4 _22020_ ( .A(_06284_ ), .Z(_07008_ ) );
BUF_X4 _22021_ ( .A(_07008_ ), .Z(_07009_ ) );
OAI22_X1 _22022_ ( .A1(_07009_ ), .A2(_05731_ ), .B1(_09105_ ), .B2(_09078_ ), .ZN(_07010_ ) );
AND3_X1 _22023_ ( .A1(_10429_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06187_ ), .ZN(_07011_ ) );
AOI221_X4 _22024_ ( .A(_07011_ ), .B1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06189_ ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06190_ ), .ZN(_07012_ ) );
NAND3_X1 _22025_ ( .A1(_06625_ ), .A2(_06460_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07013_ ) );
AOI21_X1 _22026_ ( .A(_06973_ ), .B1(_07012_ ), .B2(_07013_ ), .ZN(_07014_ ) );
AND3_X1 _22027_ ( .A1(_09068_ ), .A2(_06391_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07015_ ) );
AOI221_X4 _22028_ ( .A(_07015_ ), .B1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B2(_09122_ ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06559_ ), .ZN(_07016_ ) );
NAND3_X1 _22029_ ( .A1(_06398_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06401_ ), .ZN(_07017_ ) );
AOI21_X1 _22030_ ( .A(_06495_ ), .B1(_07016_ ), .B2(_07017_ ), .ZN(_07018_ ) );
NOR3_X1 _22031_ ( .A1(_07014_ ), .A2(_09482_ ), .A3(_07018_ ), .ZN(_07019_ ) );
NAND3_X1 _22032_ ( .A1(_06159_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06187_ ), .ZN(_07020_ ) );
INV_X1 _22033_ ( .A(_07020_ ), .ZN(_07021_ ) );
AOI221_X4 _22034_ ( .A(_07021_ ), .B1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B2(_09122_ ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06163_ ), .ZN(_07022_ ) );
NAND3_X1 _22035_ ( .A1(_06166_ ), .A2(_06167_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07023_ ) );
AOI21_X1 _22036_ ( .A(_06197_ ), .B1(_07022_ ), .B2(_07023_ ), .ZN(_07024_ ) );
AOI22_X1 _22037_ ( .A1(_06304_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06179_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07025_ ) );
AOI22_X1 _22038_ ( .A1(_06181_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_09529_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07026_ ) );
AOI21_X1 _22039_ ( .A(_06244_ ), .B1(_07025_ ), .B2(_07026_ ), .ZN(_07027_ ) );
NOR3_X1 _22040_ ( .A1(_07024_ ), .A2(_09550_ ), .A3(_07027_ ), .ZN(_07028_ ) );
NOR3_X1 _22041_ ( .A1(_07019_ ), .A2(_07028_ ), .A3(_06413_ ), .ZN(_07029_ ) );
AOI22_X1 _22042_ ( .A1(_06207_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06288_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07030_ ) );
BUF_X4 _22043_ ( .A(_09119_ ), .Z(_07031_ ) );
OAI211_X1 _22044_ ( .A(_06393_ ), .B(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06394_ ), .C2(_06395_ ), .ZN(_07032_ ) );
NAND3_X1 _22045_ ( .A1(_06407_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06408_ ), .ZN(_07033_ ) );
NAND4_X1 _22046_ ( .A1(_07030_ ), .A2(_07031_ ), .A3(_07032_ ), .A4(_07033_ ), .ZN(_07034_ ) );
AOI22_X1 _22047_ ( .A1(_06343_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06422_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07035_ ) );
AOI22_X1 _22048_ ( .A1(_06522_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06524_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07036_ ) );
NAND3_X1 _22049_ ( .A1(_07035_ ), .A2(_07036_ ), .A3(_06636_ ), .ZN(_07037_ ) );
NAND3_X1 _22050_ ( .A1(_06414_ ), .A2(_07034_ ), .A3(_07037_ ), .ZN(_07038_ ) );
AOI22_X1 _22051_ ( .A1(_06429_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06431_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07039_ ) );
OAI211_X1 _22052_ ( .A(_09094_ ), .B(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06417_ ), .C2(_06418_ ), .ZN(_07040_ ) );
NAND3_X1 _22053_ ( .A1(_06435_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06437_ ), .ZN(_07041_ ) );
NAND4_X1 _22054_ ( .A1(_07039_ ), .A2(_06433_ ), .A3(_07040_ ), .A4(_07041_ ), .ZN(_07042_ ) );
AOI22_X1 _22055_ ( .A1(_06540_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06431_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07043_ ) );
OAI211_X1 _22056_ ( .A(_09094_ ), .B(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06417_ ), .C2(_06418_ ), .ZN(_07044_ ) );
NAND3_X1 _22057_ ( .A1(_06435_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06544_ ), .ZN(_07045_ ) );
NAND4_X1 _22058_ ( .A1(_07043_ ), .A2(_06197_ ), .A3(_07044_ ), .A4(_07045_ ), .ZN(_07046_ ) );
NAND3_X1 _22059_ ( .A1(_06500_ ), .A2(_07042_ ), .A3(_07046_ ), .ZN(_07047_ ) );
AOI21_X1 _22060_ ( .A(_10252_ ), .B1(_07038_ ), .B2(_07047_ ), .ZN(_07048_ ) );
NOR3_X1 _22061_ ( .A1(_07029_ ), .A2(_06338_ ), .A3(_07048_ ), .ZN(_07049_ ) );
AND3_X1 _22062_ ( .A1(_10429_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_05809_ ), .ZN(_07050_ ) );
AOI221_X4 _22063_ ( .A(_07050_ ), .B1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_09528_ ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_09554_ ), .ZN(_07051_ ) );
NAND3_X1 _22064_ ( .A1(_06492_ ), .A2(_06167_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07052_ ) );
NAND3_X1 _22065_ ( .A1(_07051_ ), .A2(_06405_ ), .A3(_07052_ ), .ZN(_07053_ ) );
MUX2_X1 _22066_ ( .A(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .S(_06247_ ), .Z(_07054_ ) );
MUX2_X1 _22067_ ( .A(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .S(_06247_ ), .Z(_07055_ ) );
MUX2_X1 _22068_ ( .A(_07054_ ), .B(_07055_ ), .S(_10431_ ), .Z(_07056_ ) );
OAI211_X1 _22069_ ( .A(_07053_ ), .B(_09550_ ), .C1(_09085_ ), .C2(_07056_ ), .ZN(_07057_ ) );
AOI22_X1 _22070_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06522_ ), .B1(_06384_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07058_ ) );
AOI22_X1 _22071_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06638_ ), .B1(_06524_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07059_ ) );
NAND3_X1 _22072_ ( .A1(_07058_ ), .A2(_06929_ ), .A3(_07059_ ), .ZN(_07060_ ) );
BUF_X4 _22073_ ( .A(_06266_ ), .Z(_07061_ ) );
BUF_X4 _22074_ ( .A(_06383_ ), .Z(_07062_ ) );
AOI22_X1 _22075_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_07061_ ), .B1(_07062_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07063_ ) );
AOI22_X1 _22076_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06914_ ), .B1(_06915_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07064_ ) );
NAND3_X1 _22077_ ( .A1(_07063_ ), .A2(_06950_ ), .A3(_07064_ ), .ZN(_07065_ ) );
NAND3_X1 _22078_ ( .A1(_06414_ ), .A2(_07060_ ), .A3(_07065_ ), .ZN(_07066_ ) );
AOI21_X1 _22079_ ( .A(_10252_ ), .B1(_07057_ ), .B2(_07066_ ), .ZN(_07067_ ) );
AOI22_X1 _22080_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06177_ ), .B1(_06504_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07068_ ) );
AOI22_X1 _22081_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06288_ ), .B1(_06506_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07069_ ) );
AOI21_X1 _22082_ ( .A(_06284_ ), .B1(_07068_ ), .B2(_07069_ ), .ZN(_07070_ ) );
AOI22_X1 _22083_ ( .A1(_06177_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06179_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07071_ ) );
AOI22_X1 _22084_ ( .A1(_06181_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_09529_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07072_ ) );
AOI21_X1 _22085_ ( .A(_09084_ ), .B1(_07071_ ), .B2(_07072_ ), .ZN(_07073_ ) );
OAI21_X1 _22086_ ( .A(_09482_ ), .B1(_07070_ ), .B2(_07073_ ), .ZN(_07074_ ) );
AOI22_X1 _22087_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06304_ ), .B1(_06504_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07075_ ) );
AOI22_X1 _22088_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06179_ ), .B1(_09529_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07076_ ) );
AOI21_X1 _22089_ ( .A(_09084_ ), .B1(_07075_ ), .B2(_07076_ ), .ZN(_07077_ ) );
AOI22_X1 _22090_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06304_ ), .B1(_06504_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07078_ ) );
AOI22_X1 _22091_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06179_ ), .B1(_09529_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07079_ ) );
AOI21_X1 _22092_ ( .A(_06244_ ), .B1(_07078_ ), .B2(_07079_ ), .ZN(_07080_ ) );
OAI21_X1 _22093_ ( .A(_09550_ ), .B1(_07077_ ), .B2(_07080_ ), .ZN(_07081_ ) );
AOI21_X1 _22094_ ( .A(_09664_ ), .B1(_07074_ ), .B2(_07081_ ), .ZN(_07082_ ) );
NOR3_X1 _22095_ ( .A1(_07067_ ), .A2(_07082_ ), .A3(_10009_ ), .ZN(_07083_ ) );
NOR3_X1 _22096_ ( .A1(_07049_ ), .A2(_07083_ ), .A3(_09020_ ), .ZN(_07084_ ) );
AND3_X1 _22097_ ( .A1(_06228_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06229_ ), .ZN(_07085_ ) );
AOI221_X4 _22098_ ( .A(_07085_ ), .B1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06231_ ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06285_ ), .ZN(_07086_ ) );
NAND3_X1 _22099_ ( .A1(_06568_ ), .A2(_06236_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07087_ ) );
NAND3_X1 _22100_ ( .A1(_07086_ ), .A2(_06611_ ), .A3(_07087_ ), .ZN(_07088_ ) );
AND3_X1 _22101_ ( .A1(_06456_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06240_ ), .ZN(_07089_ ) );
AOI221_X4 _22102_ ( .A(_07089_ ), .B1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06923_ ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06176_ ), .ZN(_07090_ ) );
NAND3_X1 _22103_ ( .A1(_06925_ ), .A2(_06811_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07091_ ) );
NAND3_X1 _22104_ ( .A1(_07090_ ), .A2(_06596_ ), .A3(_07091_ ), .ZN(_07092_ ) );
NAND3_X1 _22105_ ( .A1(_07088_ ), .A2(_07092_ ), .A3(_06684_ ), .ZN(_07093_ ) );
AOI22_X1 _22106_ ( .A1(_06836_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_09484_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07094_ ) );
OAI211_X1 _22107_ ( .A(_06978_ ), .B(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06394_ ), .C2(_06395_ ), .ZN(_07095_ ) );
NAND3_X1 _22108_ ( .A1(_06492_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06931_ ), .ZN(_07096_ ) );
NAND4_X1 _22109_ ( .A1(_07094_ ), .A2(_06973_ ), .A3(_07095_ ), .A4(_07096_ ), .ZN(_07097_ ) );
AOI22_X1 _22110_ ( .A1(_06342_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06470_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07098_ ) );
AOI22_X1 _22111_ ( .A1(_06609_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06213_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07099_ ) );
NAND3_X1 _22112_ ( .A1(_07098_ ), .A2(_07099_ ), .A3(_06964_ ), .ZN(_07100_ ) );
NAND3_X1 _22113_ ( .A1(_06254_ ), .A2(_07097_ ), .A3(_07100_ ), .ZN(_07101_ ) );
AOI21_X1 _22114_ ( .A(_09665_ ), .B1(_07093_ ), .B2(_07101_ ), .ZN(_07102_ ) );
AOI22_X1 _22115_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06216_ ), .B1(_06649_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07103_ ) );
AOI22_X1 _22116_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06220_ ), .B1(_06221_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07104_ ) );
NAND3_X1 _22117_ ( .A1(_07103_ ), .A2(_06479_ ), .A3(_07104_ ), .ZN(_07105_ ) );
AOI22_X1 _22118_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06369_ ), .B1(_06702_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07106_ ) );
AOI22_X1 _22119_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_07061_ ), .B1(_07062_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07107_ ) );
NAND3_X1 _22120_ ( .A1(_07106_ ), .A2(_06192_ ), .A3(_07107_ ), .ZN(_07108_ ) );
NAND3_X1 _22121_ ( .A1(_06254_ ), .A2(_07105_ ), .A3(_07108_ ), .ZN(_07109_ ) );
AOI22_X1 _22122_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06220_ ), .B1(_06221_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07110_ ) );
AOI22_X1 _22123_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06444_ ), .B1(_06527_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07111_ ) );
NAND3_X1 _22124_ ( .A1(_07110_ ), .A2(_06514_ ), .A3(_07111_ ), .ZN(_07112_ ) );
AOI22_X1 _22125_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06522_ ), .B1(_07062_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07113_ ) );
AOI22_X1 _22126_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06638_ ), .B1(_06524_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07114_ ) );
NAND3_X1 _22127_ ( .A1(_07113_ ), .A2(_06950_ ), .A3(_07114_ ), .ZN(_07115_ ) );
NAND3_X1 _22128_ ( .A1(_06388_ ), .A2(_07112_ ), .A3(_07115_ ), .ZN(_07116_ ) );
AOI21_X1 _22129_ ( .A(_10252_ ), .B1(_07109_ ), .B2(_07116_ ), .ZN(_07117_ ) );
OAI21_X1 _22130_ ( .A(_06227_ ), .B1(_07102_ ), .B2(_07117_ ), .ZN(_07118_ ) );
AOI22_X1 _22131_ ( .A1(_06836_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_09484_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07119_ ) );
OAI211_X1 _22132_ ( .A(_06939_ ), .B(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06480_ ), .C2(_06481_ ), .ZN(_07120_ ) );
NAND3_X1 _22133_ ( .A1(_06492_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06931_ ), .ZN(_07121_ ) );
NAND4_X1 _22134_ ( .A1(_07119_ ), .A2(_06973_ ), .A3(_07120_ ), .A4(_07121_ ), .ZN(_07122_ ) );
AOI22_X1 _22135_ ( .A1(_06836_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06422_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07123_ ) );
OAI211_X1 _22136_ ( .A(_06978_ ), .B(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06394_ ), .C2(_06395_ ), .ZN(_07124_ ) );
NAND3_X1 _22137_ ( .A1(_06398_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06931_ ), .ZN(_07125_ ) );
NAND4_X1 _22138_ ( .A1(_07123_ ), .A2(_06255_ ), .A3(_07124_ ), .A4(_07125_ ), .ZN(_07126_ ) );
NAND3_X1 _22139_ ( .A1(_06254_ ), .A2(_07122_ ), .A3(_07126_ ), .ZN(_07127_ ) );
AOI22_X1 _22140_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06794_ ), .B1(_06274_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07128_ ) );
AOI22_X1 _22141_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06267_ ), .B1(_09795_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07129_ ) );
NAND3_X1 _22142_ ( .A1(_07128_ ), .A2(_06144_ ), .A3(_07129_ ), .ZN(_07130_ ) );
AOI22_X1 _22143_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06382_ ), .B1(_06540_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07131_ ) );
AOI22_X1 _22144_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06477_ ), .B1(_06425_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07132_ ) );
NAND3_X1 _22145_ ( .A1(_07131_ ), .A2(_06700_ ), .A3(_07132_ ), .ZN(_07133_ ) );
NAND3_X1 _22146_ ( .A1(_06388_ ), .A2(_07130_ ), .A3(_07133_ ), .ZN(_07134_ ) );
AOI21_X1 _22147_ ( .A(_06186_ ), .B1(_07127_ ), .B2(_07134_ ), .ZN(_07135_ ) );
AOI22_X1 _22148_ ( .A1(_06522_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06524_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07136_ ) );
NAND3_X1 _22149_ ( .A1(_06407_ ), .A2(_06939_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07137_ ) );
NAND3_X1 _22150_ ( .A1(_06441_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06408_ ), .ZN(_07138_ ) );
NAND4_X1 _22151_ ( .A1(_07136_ ), .A2(_06390_ ), .A3(_07137_ ), .A4(_07138_ ), .ZN(_07139_ ) );
AOI22_X1 _22152_ ( .A1(_07061_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06915_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07140_ ) );
NAND3_X1 _22153_ ( .A1(_06441_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06408_ ), .ZN(_07141_ ) );
NAND3_X1 _22154_ ( .A1(_06407_ ), .A2(_06978_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07142_ ) );
NAND4_X1 _22155_ ( .A1(_07140_ ), .A2(_07031_ ), .A3(_07141_ ), .A4(_07142_ ), .ZN(_07143_ ) );
NAND3_X1 _22156_ ( .A1(_06414_ ), .A2(_07139_ ), .A3(_07143_ ), .ZN(_07144_ ) );
AOI22_X1 _22157_ ( .A1(_06444_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06431_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07145_ ) );
OAI211_X1 _22158_ ( .A(_09094_ ), .B(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06417_ ), .C2(_06418_ ), .ZN(_07146_ ) );
NAND3_X1 _22159_ ( .A1(_06435_ ), .A2(_06393_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07147_ ) );
NAND4_X1 _22160_ ( .A1(_07145_ ), .A2(_06433_ ), .A3(_07146_ ), .A4(_07147_ ), .ZN(_07148_ ) );
AOI22_X1 _22161_ ( .A1(_06522_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06288_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07149_ ) );
AOI22_X1 _22162_ ( .A1(_06649_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06445_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07150_ ) );
NAND3_X1 _22163_ ( .A1(_07149_ ), .A2(_07150_ ), .A3(_07031_ ), .ZN(_07151_ ) );
NAND3_X1 _22164_ ( .A1(_09463_ ), .A2(_07148_ ), .A3(_07151_ ), .ZN(_07152_ ) );
AOI21_X1 _22165_ ( .A(_06413_ ), .B1(_07144_ ), .B2(_07152_ ), .ZN(_07153_ ) );
OAI21_X1 _22166_ ( .A(_06338_ ), .B1(_07135_ ), .B2(_07153_ ), .ZN(_07154_ ) );
AOI21_X1 _22167_ ( .A(_09604_ ), .B1(_07118_ ), .B2(_07154_ ), .ZN(_07155_ ) );
OAI21_X1 _22168_ ( .A(_09138_ ), .B1(_07084_ ), .B2(_07155_ ), .ZN(_07156_ ) );
AND3_X1 _22169_ ( .A1(_06456_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06240_ ), .ZN(_07157_ ) );
AOI221_X4 _22170_ ( .A(_07157_ ), .B1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06923_ ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06176_ ), .ZN(_07158_ ) );
NAND3_X1 _22171_ ( .A1(_06925_ ), .A2(_06811_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07159_ ) );
NAND3_X1 _22172_ ( .A1(_07158_ ), .A2(_06308_ ), .A3(_07159_ ), .ZN(_07160_ ) );
MUX2_X1 _22173_ ( .A(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .S(_06464_ ), .Z(_07161_ ) );
MUX2_X1 _22174_ ( .A(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .S(_06464_ ), .Z(_07162_ ) );
MUX2_X1 _22175_ ( .A(_07161_ ), .B(_07162_ ), .S(_06448_ ), .Z(_07163_ ) );
OAI211_X1 _22176_ ( .A(_07160_ ), .B(_06252_ ), .C1(_06198_ ), .C2(_07163_ ), .ZN(_07164_ ) );
NAND3_X1 _22177_ ( .A1(_06145_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06146_ ), .ZN(_07165_ ) );
INV_X1 _22178_ ( .A(_07165_ ), .ZN(_07166_ ) );
AOI221_X4 _22179_ ( .A(_07166_ ), .B1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06149_ ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06424_ ), .ZN(_07167_ ) );
NAND3_X1 _22180_ ( .A1(_06925_ ), .A2(_06811_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07168_ ) );
AOI21_X1 _22181_ ( .A(_06479_ ), .B1(_07167_ ), .B2(_07168_ ), .ZN(_07169_ ) );
OAI211_X1 _22182_ ( .A(_06160_ ), .B(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06629_ ), .C2(_06630_ ), .ZN(_07170_ ) );
INV_X1 _22183_ ( .A(_07170_ ), .ZN(_07171_ ) );
AOI221_X4 _22184_ ( .A(_07171_ ), .B1(_06923_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C2(_09626_ ), .ZN(_07172_ ) );
NAND3_X1 _22185_ ( .A1(_06330_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06783_ ), .ZN(_07173_ ) );
AOI21_X1 _22186_ ( .A(_06255_ ), .B1(_07172_ ), .B2(_07173_ ), .ZN(_07174_ ) );
OAI21_X1 _22187_ ( .A(_06890_ ), .B1(_07169_ ), .B2(_07174_ ), .ZN(_07175_ ) );
AOI21_X1 _22188_ ( .A(_09487_ ), .B1(_07164_ ), .B2(_07175_ ), .ZN(_07176_ ) );
NAND3_X1 _22189_ ( .A1(_06145_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06678_ ), .ZN(_07177_ ) );
INV_X1 _22190_ ( .A(_07177_ ), .ZN(_07178_ ) );
AOI221_X4 _22191_ ( .A(_07178_ ), .B1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06178_ ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06150_ ), .ZN(_07179_ ) );
NAND3_X1 _22192_ ( .A1(_06152_ ), .A2(_06460_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07180_ ) );
AOI21_X1 _22193_ ( .A(_06144_ ), .B1(_07179_ ), .B2(_07180_ ), .ZN(_07181_ ) );
NAND3_X1 _22194_ ( .A1(_06239_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06240_ ), .ZN(_07182_ ) );
INV_X1 _22195_ ( .A(_07182_ ), .ZN(_07183_ ) );
AOI221_X4 _22196_ ( .A(_07183_ ), .B1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06178_ ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06259_ ), .ZN(_07184_ ) );
NAND3_X1 _22197_ ( .A1(_06193_ ), .A2(_06194_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07185_ ) );
AOI21_X1 _22198_ ( .A(_06390_ ), .B1(_07184_ ), .B2(_07185_ ), .ZN(_07186_ ) );
OAI21_X1 _22199_ ( .A(_06645_ ), .B1(_07181_ ), .B2(_07186_ ), .ZN(_07187_ ) );
AOI22_X1 _22200_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06421_ ), .B1(_06649_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07188_ ) );
AOI22_X1 _22201_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06347_ ), .B1(_06640_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07189_ ) );
AOI21_X1 _22202_ ( .A(_06255_ ), .B1(_07188_ ), .B2(_07189_ ), .ZN(_07190_ ) );
AOI22_X1 _22203_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_07061_ ), .B1(_09795_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07191_ ) );
AOI22_X1 _22204_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06914_ ), .B1(_06915_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07192_ ) );
AOI21_X1 _22205_ ( .A(_06158_ ), .B1(_07191_ ), .B2(_07192_ ), .ZN(_07193_ ) );
OAI21_X1 _22206_ ( .A(_06684_ ), .B1(_07190_ ), .B2(_07193_ ), .ZN(_07194_ ) );
AOI21_X1 _22207_ ( .A(_09665_ ), .B1(_07187_ ), .B2(_07194_ ), .ZN(_07195_ ) );
OAI21_X1 _22208_ ( .A(_06143_ ), .B1(_07176_ ), .B2(_07195_ ), .ZN(_07196_ ) );
AND3_X1 _22209_ ( .A1(_06557_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06146_ ), .ZN(_07197_ ) );
AOI221_X4 _22210_ ( .A(_07197_ ), .B1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06716_ ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06266_ ), .ZN(_07198_ ) );
NAND3_X1 _22211_ ( .A1(_06718_ ), .A2(_06562_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07199_ ) );
AOI21_X1 _22212_ ( .A(_06245_ ), .B1(_07198_ ), .B2(_07199_ ), .ZN(_07200_ ) );
AND3_X1 _22213_ ( .A1(_06239_ ), .A2(_06391_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07201_ ) );
AOI221_X4 _22214_ ( .A(_07201_ ), .B1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06149_ ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06424_ ), .ZN(_07202_ ) );
NAND3_X1 _22215_ ( .A1(_06568_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06736_ ), .ZN(_07203_ ) );
AOI21_X1 _22216_ ( .A(_06329_ ), .B1(_07202_ ), .B2(_07203_ ), .ZN(_07204_ ) );
OAI21_X1 _22217_ ( .A(_06555_ ), .B1(_07200_ ), .B2(_07204_ ), .ZN(_07205_ ) );
OAI211_X1 _22218_ ( .A(_06678_ ), .B(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06351_ ), .C2(_06354_ ), .ZN(_07206_ ) );
INV_X1 _22219_ ( .A(_07206_ ), .ZN(_07207_ ) );
AOI221_X4 _22220_ ( .A(_07207_ ), .B1(_06716_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06285_ ), .ZN(_07208_ ) );
NAND3_X1 _22221_ ( .A1(_06235_ ), .A2(_06236_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07209_ ) );
AOI21_X1 _22222_ ( .A(_06565_ ), .B1(_07208_ ), .B2(_07209_ ), .ZN(_07210_ ) );
AOI22_X1 _22223_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06365_ ), .B1(_06366_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07211_ ) );
AOI22_X1 _22224_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06594_ ), .B1(_06370_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07212_ ) );
AOI21_X1 _22225_ ( .A(_06144_ ), .B1(_07211_ ), .B2(_07212_ ), .ZN(_07213_ ) );
OAI21_X1 _22226_ ( .A(_06573_ ), .B1(_07210_ ), .B2(_07213_ ), .ZN(_07214_ ) );
NAND3_X1 _22227_ ( .A1(_07205_ ), .A2(_09784_ ), .A3(_07214_ ), .ZN(_07215_ ) );
NAND3_X1 _22228_ ( .A1(_06671_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06399_ ), .ZN(_07216_ ) );
INV_X1 _22229_ ( .A(_07216_ ), .ZN(_07217_ ) );
AOI221_X4 _22230_ ( .A(_07217_ ), .B1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06430_ ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06326_ ), .ZN(_07218_ ) );
NAND3_X1 _22231_ ( .A1(_09071_ ), .A2(_09095_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07219_ ) );
NAND3_X1 _22232_ ( .A1(_07218_ ), .A2(_09085_ ), .A3(_07219_ ), .ZN(_07220_ ) );
NAND3_X1 _22233_ ( .A1(_06671_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06399_ ), .ZN(_07221_ ) );
INV_X1 _22234_ ( .A(_07221_ ), .ZN(_07222_ ) );
AOI221_X4 _22235_ ( .A(_07222_ ), .B1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06430_ ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06326_ ), .ZN(_07223_ ) );
NAND3_X1 _22236_ ( .A1(_06561_ ), .A2(_06562_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07224_ ) );
NAND3_X1 _22237_ ( .A1(_07223_ ), .A2(_06300_ ), .A3(_07224_ ), .ZN(_07225_ ) );
NAND3_X1 _22238_ ( .A1(_07220_ ), .A2(_07225_ ), .A3(_06303_ ), .ZN(_07226_ ) );
AOI22_X1 _22239_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06342_ ), .B1(_06263_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07227_ ) );
AOI22_X1 _22240_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06379_ ), .B1(_06380_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07228_ ) );
AOI21_X1 _22241_ ( .A(_06192_ ), .B1(_07227_ ), .B2(_07228_ ), .ZN(_07229_ ) );
AOI22_X1 _22242_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06421_ ), .B1(_06649_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07230_ ) );
AOI22_X1 _22243_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06347_ ), .B1(_06640_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07231_ ) );
AOI21_X1 _22244_ ( .A(_06636_ ), .B1(_07230_ ), .B2(_07231_ ), .ZN(_07232_ ) );
OAI21_X1 _22245_ ( .A(_06890_ ), .B1(_07229_ ), .B2(_07232_ ), .ZN(_07233_ ) );
NAND3_X1 _22246_ ( .A1(_07226_ ), .A2(_11056_ ), .A3(_07233_ ), .ZN(_07234_ ) );
NAND3_X1 _22247_ ( .A1(_07215_ ), .A2(_10744_ ), .A3(_07234_ ), .ZN(_07235_ ) );
NAND3_X1 _22248_ ( .A1(_07196_ ), .A2(_07235_ ), .A3(_02457_ ), .ZN(_07236_ ) );
AND3_X1 _22249_ ( .A1(_10429_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06187_ ), .ZN(_07237_ ) );
AOI221_X4 _22250_ ( .A(_07237_ ), .B1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06189_ ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06190_ ), .ZN(_07238_ ) );
NAND3_X1 _22251_ ( .A1(_06330_ ), .A2(_06331_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07239_ ) );
NAND3_X1 _22252_ ( .A1(_07238_ ), .A2(_06964_ ), .A3(_07239_ ), .ZN(_07240_ ) );
MUX2_X1 _22253_ ( .A(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .S(_06199_ ), .Z(_07241_ ) );
MUX2_X1 _22254_ ( .A(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .S(_06199_ ), .Z(_07242_ ) );
MUX2_X1 _22255_ ( .A(_07241_ ), .B(_07242_ ), .S(_06448_ ), .Z(_07243_ ) );
OAI211_X1 _22256_ ( .A(_07240_ ), .B(_06414_ ), .C1(_06198_ ), .C2(_07243_ ), .ZN(_07244_ ) );
AOI22_X1 _22257_ ( .A1(_06232_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06259_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07245_ ) );
NAND3_X1 _22258_ ( .A1(_06440_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06400_ ), .ZN(_07246_ ) );
NAND3_X1 _22259_ ( .A1(_06397_ ), .A2(_06598_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07247_ ) );
AND3_X1 _22260_ ( .A1(_07245_ ), .A2(_07246_ ), .A3(_07247_ ), .ZN(_07248_ ) );
AOI22_X1 _22261_ ( .A1(_06266_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06150_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07249_ ) );
NAND3_X1 _22262_ ( .A1(_06440_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06400_ ), .ZN(_07250_ ) );
NAND3_X1 _22263_ ( .A1(_06397_ ), .A2(_06598_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07251_ ) );
AND3_X1 _22264_ ( .A1(_07249_ ), .A2(_07250_ ), .A3(_07251_ ), .ZN(_07252_ ) );
MUX2_X1 _22265_ ( .A(_07248_ ), .B(_07252_ ), .S(_06433_ ), .Z(_07253_ ) );
OAI211_X1 _22266_ ( .A(_07244_ ), .B(_06654_ ), .C1(_10529_ ), .C2(_07253_ ), .ZN(_07254_ ) );
AND3_X1 _22267_ ( .A1(_06228_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06229_ ), .ZN(_07255_ ) );
AOI221_X4 _22268_ ( .A(_07255_ ), .B1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06231_ ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06232_ ), .ZN(_07256_ ) );
NAND3_X1 _22269_ ( .A1(_06235_ ), .A2(_06236_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07257_ ) );
AOI21_X1 _22270_ ( .A(_06362_ ), .B1(_07256_ ), .B2(_07257_ ), .ZN(_07258_ ) );
AND3_X1 _22271_ ( .A1(_06456_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06240_ ), .ZN(_07259_ ) );
AOI221_X4 _22272_ ( .A(_07259_ ), .B1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06923_ ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06176_ ), .ZN(_07260_ ) );
NAND3_X1 _22273_ ( .A1(_06309_ ), .A2(_06154_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07261_ ) );
AOI21_X1 _22274_ ( .A(_06479_ ), .B1(_07260_ ), .B2(_07261_ ), .ZN(_07262_ ) );
OAI21_X1 _22275_ ( .A(_06555_ ), .B1(_07258_ ), .B2(_07262_ ), .ZN(_07263_ ) );
AND3_X1 _22276_ ( .A1(_06456_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06160_ ), .ZN(_07264_ ) );
AOI221_X4 _22277_ ( .A(_07264_ ), .B1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06189_ ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06190_ ), .ZN(_07265_ ) );
NAND3_X1 _22278_ ( .A1(_06459_ ), .A2(_06460_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07266_ ) );
NAND3_X1 _22279_ ( .A1(_07265_ ), .A2(_06362_ ), .A3(_07266_ ), .ZN(_07267_ ) );
AOI22_X1 _22280_ ( .A1(_06205_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06274_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07268_ ) );
OAI211_X1 _22281_ ( .A(_06798_ ), .B(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06353_ ), .C2(_06356_ ), .ZN(_07269_ ) );
NAND3_X1 _22282_ ( .A1(_06193_ ), .A2(_06194_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07270_ ) );
NAND3_X1 _22283_ ( .A1(_07268_ ), .A2(_07269_ ), .A3(_07270_ ), .ZN(_07271_ ) );
OAI211_X1 _22284_ ( .A(_07267_ ), .B(_06463_ ), .C1(_06198_ ), .C2(_07271_ ), .ZN(_07272_ ) );
NAND3_X1 _22285_ ( .A1(_07263_ ), .A2(_10053_ ), .A3(_07272_ ), .ZN(_07273_ ) );
NAND3_X1 _22286_ ( .A1(_07254_ ), .A2(_07273_ ), .A3(_06143_ ), .ZN(_07274_ ) );
NAND3_X1 _22287_ ( .A1(_06239_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06229_ ), .ZN(_07275_ ) );
INV_X1 _22288_ ( .A(_07275_ ), .ZN(_07276_ ) );
AOI221_X4 _22289_ ( .A(_07276_ ), .B1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06178_ ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06259_ ), .ZN(_07277_ ) );
NAND3_X1 _22290_ ( .A1(_06625_ ), .A2(_06331_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07278_ ) );
AOI21_X1 _22291_ ( .A(_06950_ ), .B1(_07277_ ), .B2(_07278_ ), .ZN(_07279_ ) );
NAND3_X1 _22292_ ( .A1(_06159_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06240_ ), .ZN(_07280_ ) );
INV_X1 _22293_ ( .A(_07280_ ), .ZN(_07281_ ) );
AOI221_X4 _22294_ ( .A(_07281_ ), .B1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06178_ ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06259_ ), .ZN(_07282_ ) );
NAND3_X1 _22295_ ( .A1(_06483_ ), .A2(_06599_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07283_ ) );
AOI21_X1 _22296_ ( .A(_07031_ ), .B1(_07282_ ), .B2(_07283_ ), .ZN(_07284_ ) );
OAI21_X1 _22297_ ( .A(_06204_ ), .B1(_07279_ ), .B2(_07284_ ), .ZN(_07285_ ) );
AND3_X1 _22298_ ( .A1(_06159_ ), .A2(_06391_ ), .A3(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07286_ ) );
AOI221_X4 _22299_ ( .A(_07286_ ), .B1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_09528_ ), .C1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06190_ ), .ZN(_07287_ ) );
NAND3_X1 _22300_ ( .A1(_06725_ ), .A2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06798_ ), .ZN(_07288_ ) );
NAND3_X1 _22301_ ( .A1(_07287_ ), .A2(_06929_ ), .A3(_07288_ ), .ZN(_07289_ ) );
MUX2_X1 _22302_ ( .A(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .S(_06247_ ), .Z(_07290_ ) );
MUX2_X1 _22303_ ( .A(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .S(_06247_ ), .Z(_07291_ ) );
MUX2_X1 _22304_ ( .A(_07290_ ), .B(_07291_ ), .S(_10431_ ), .Z(_07292_ ) );
OAI211_X1 _22305_ ( .A(_07289_ ), .B(_06500_ ), .C1(_09085_ ), .C2(_07292_ ), .ZN(_07293_ ) );
AOI21_X1 _22306_ ( .A(_09665_ ), .B1(_07285_ ), .B2(_07293_ ), .ZN(_07294_ ) );
AOI22_X1 _22307_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06522_ ), .B1(_07062_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07295_ ) );
AOI22_X1 _22308_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06638_ ), .B1(_06524_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07296_ ) );
AOI21_X1 _22309_ ( .A(_07031_ ), .B1(_07295_ ), .B2(_07296_ ), .ZN(_07297_ ) );
AOI22_X1 _22310_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06286_ ), .B1(_06527_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07298_ ) );
AOI22_X1 _22311_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06422_ ), .B1(_06445_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07299_ ) );
AOI21_X1 _22312_ ( .A(_06284_ ), .B1(_07298_ ), .B2(_07299_ ), .ZN(_07300_ ) );
OAI21_X1 _22313_ ( .A(_06414_ ), .B1(_07297_ ), .B2(_07300_ ), .ZN(_07301_ ) );
AOI22_X1 _22314_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06382_ ), .B1(_06384_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07302_ ) );
AOI22_X1 _22315_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06477_ ), .B1(_06524_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07303_ ) );
NAND3_X1 _22316_ ( .A1(_07302_ ), .A2(_06973_ ), .A3(_07303_ ), .ZN(_07304_ ) );
AOI22_X1 _22317_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06522_ ), .B1(_07062_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07305_ ) );
AOI22_X1 _22318_ ( .A1(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06638_ ), .B1(_06915_ ), .B2(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07306_ ) );
NAND3_X1 _22319_ ( .A1(_07305_ ), .A2(_06929_ ), .A3(_07306_ ), .ZN(_07307_ ) );
NAND3_X1 _22320_ ( .A1(_06388_ ), .A2(_07304_ ), .A3(_07307_ ), .ZN(_07308_ ) );
AOI21_X1 _22321_ ( .A(_10252_ ), .B1(_07301_ ), .B2(_07308_ ), .ZN(_07309_ ) );
OAI21_X1 _22322_ ( .A(_06227_ ), .B1(_07294_ ), .B2(_07309_ ), .ZN(_07310_ ) );
NAND3_X1 _22323_ ( .A1(_07274_ ), .A2(_09604_ ), .A3(_07310_ ), .ZN(_07311_ ) );
NAND3_X1 _22324_ ( .A1(_07236_ ), .A2(_07311_ ), .A3(_09035_ ), .ZN(_07312_ ) );
AND3_X1 _22325_ ( .A1(_07156_ ), .A2(_06077_ ), .A3(_07312_ ), .ZN(\load_data_out[4] ) );
INV_X1 _22326_ ( .A(\load_data_out[4] ), .ZN(_07313_ ) );
OAI21_X1 _22327_ ( .A(_07313_ ), .B1(_07009_ ), .B2(_06130_ ), .ZN(_07314_ ) );
AOI21_X1 _22328_ ( .A(_07010_ ), .B1(_07314_ ), .B2(_06102_ ), .ZN(_07315_ ) );
NOR2_X1 _22329_ ( .A1(_07315_ ), .A2(_06137_ ), .ZN(_00025_ ) );
OAI22_X1 _22330_ ( .A1(_10433_ ), .A2(_05731_ ), .B1(_09105_ ), .B2(_09074_ ), .ZN(_07316_ ) );
AND3_X1 _22331_ ( .A1(_06557_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06678_ ), .ZN(_07317_ ) );
AOI221_X4 _22332_ ( .A(_07317_ ), .B1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06559_ ), .C1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06232_ ), .ZN(_07318_ ) );
NAND3_X1 _22333_ ( .A1(_06561_ ), .A2(_06562_ ), .A3(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07319_ ) );
AOI21_X1 _22334_ ( .A(_06362_ ), .B1(_07318_ ), .B2(_07319_ ), .ZN(_07320_ ) );
AND3_X1 _22335_ ( .A1(_10429_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06187_ ), .ZN(_07321_ ) );
AOI221_X4 _22336_ ( .A(_07321_ ), .B1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06189_ ), .C1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06190_ ), .ZN(_07322_ ) );
NAND3_X1 _22337_ ( .A1(_06625_ ), .A2(_06460_ ), .A3(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07323_ ) );
AOI21_X1 _22338_ ( .A(_06973_ ), .B1(_07322_ ), .B2(_07323_ ), .ZN(_07324_ ) );
NOR3_X1 _22339_ ( .A1(_07320_ ), .A2(_07324_ ), .A3(_06463_ ), .ZN(_07325_ ) );
NAND3_X1 _22340_ ( .A1(_06239_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06256_ ), .ZN(_07326_ ) );
INV_X1 _22341_ ( .A(_07326_ ), .ZN(_07327_ ) );
AOI221_X4 _22342_ ( .A(_07327_ ), .B1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06178_ ), .C1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06259_ ), .ZN(_07328_ ) );
NAND3_X1 _22343_ ( .A1(_06193_ ), .A2(_06194_ ), .A3(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07329_ ) );
AOI21_X1 _22344_ ( .A(_06636_ ), .B1(_07328_ ), .B2(_07329_ ), .ZN(_07330_ ) );
NAND3_X1 _22345_ ( .A1(_06159_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06187_ ), .ZN(_07331_ ) );
INV_X1 _22346_ ( .A(_07331_ ), .ZN(_07332_ ) );
AOI221_X4 _22347_ ( .A(_07332_ ), .B1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B2(_09122_ ), .C1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06559_ ), .ZN(_07333_ ) );
NAND3_X1 _22348_ ( .A1(_06398_ ), .A2(_06350_ ), .A3(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07334_ ) );
AOI21_X1 _22349_ ( .A(_06495_ ), .B1(_07333_ ), .B2(_07334_ ), .ZN(_07335_ ) );
NOR3_X1 _22350_ ( .A1(_07330_ ), .A2(_07335_ ), .A3(_09550_ ), .ZN(_07336_ ) );
NOR3_X1 _22351_ ( .A1(_07325_ ), .A2(_06654_ ), .A3(_07336_ ), .ZN(_07337_ ) );
AOI22_X1 _22352_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06382_ ), .B1(_06540_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07338_ ) );
AOI22_X1 _22353_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06470_ ), .B1(_06864_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07339_ ) );
AOI21_X1 _22354_ ( .A(_06405_ ), .B1(_07338_ ), .B2(_07339_ ), .ZN(_07340_ ) );
AOI22_X1 _22355_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06267_ ), .B1(_09795_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07341_ ) );
AOI22_X1 _22356_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_09484_ ), .B1(_06268_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07342_ ) );
AOI21_X1 _22357_ ( .A(_06158_ ), .B1(_07341_ ), .B2(_07342_ ), .ZN(_07343_ ) );
NOR3_X1 _22358_ ( .A1(_06890_ ), .A2(_07340_ ), .A3(_07343_ ), .ZN(_07344_ ) );
AOI22_X1 _22359_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06286_ ), .B1(_06181_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07345_ ) );
AOI22_X1 _22360_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06288_ ), .B1(_06289_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07346_ ) );
AOI21_X1 _22361_ ( .A(_06495_ ), .B1(_07345_ ), .B2(_07346_ ), .ZN(_07347_ ) );
AOI22_X1 _22362_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06177_ ), .B1(_06504_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07348_ ) );
AOI22_X1 _22363_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06431_ ), .B1(_06506_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07349_ ) );
AOI21_X1 _22364_ ( .A(_06284_ ), .B1(_07348_ ), .B2(_07349_ ), .ZN(_07350_ ) );
NOR3_X1 _22365_ ( .A1(_06388_ ), .A2(_07347_ ), .A3(_07350_ ), .ZN(_07351_ ) );
NOR3_X1 _22366_ ( .A1(_07344_ ), .A2(_07351_ ), .A3(_09594_ ), .ZN(_07352_ ) );
OAI21_X1 _22367_ ( .A(_09489_ ), .B1(_07337_ ), .B2(_07352_ ), .ZN(_07353_ ) );
AOI22_X1 _22368_ ( .A1(_06316_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06306_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07354_ ) );
OAI211_X1 _22369_ ( .A(_06333_ ), .B(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06587_ ), .C2(_06588_ ), .ZN(_07355_ ) );
NAND3_X1 _22370_ ( .A1(_06625_ ), .A2(_06460_ ), .A3(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07356_ ) );
NAND4_X1 _22371_ ( .A1(_07354_ ), .A2(_06368_ ), .A3(_07355_ ), .A4(_07356_ ), .ZN(_07357_ ) );
AOI22_X1 _22372_ ( .A1(_06574_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06325_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07358_ ) );
AOI22_X1 _22373_ ( .A1(_06593_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06306_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07359_ ) );
NAND3_X1 _22374_ ( .A1(_07358_ ), .A2(_07359_ ), .A3(_06611_ ), .ZN(_07360_ ) );
NAND3_X1 _22375_ ( .A1(_06555_ ), .A2(_07357_ ), .A3(_07360_ ), .ZN(_07361_ ) );
BUF_X2 _22376_ ( .A(_10430_ ), .Z(_07362_ ) );
AND3_X1 _22377_ ( .A1(_07362_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06248_ ), .ZN(_07363_ ) );
OAI211_X1 _22378_ ( .A(_06392_ ), .B(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06352_ ), .C2(_06355_ ), .ZN(_07364_ ) );
NAND3_X1 _22379_ ( .A1(_06397_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06400_ ), .ZN(_07365_ ) );
NAND2_X1 _22380_ ( .A1(_07364_ ), .A2(_07365_ ), .ZN(_07366_ ) );
AND3_X1 _22381_ ( .A1(_06434_ ), .A2(_06392_ ), .A3(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07367_ ) );
NOR3_X1 _22382_ ( .A1(_07363_ ), .A2(_07366_ ), .A3(_07367_ ), .ZN(_07368_ ) );
AOI22_X1 _22383_ ( .A1(_09745_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06326_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07369_ ) );
NAND3_X1 _22384_ ( .A1(_06165_ ), .A2(_06153_ ), .A3(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07370_ ) );
NAND3_X1 _22385_ ( .A1(_07362_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06248_ ), .ZN(_07371_ ) );
AND3_X1 _22386_ ( .A1(_07369_ ), .A2(_07370_ ), .A3(_07371_ ), .ZN(_07372_ ) );
MUX2_X1 _22387_ ( .A(_07368_ ), .B(_07372_ ), .S(_06973_ ), .Z(_07373_ ) );
OAI211_X1 _22388_ ( .A(_10053_ ), .B(_07361_ ), .C1(_07373_ ), .C2(_09744_ ), .ZN(_07374_ ) );
AOI22_X1 _22389_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06574_ ), .B1(_06781_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07375_ ) );
AOI22_X1 _22390_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06339_ ), .B1(_09530_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07376_ ) );
AOI21_X1 _22391_ ( .A(_06611_ ), .B1(_07375_ ), .B2(_07376_ ), .ZN(_07377_ ) );
AOI22_X1 _22392_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06605_ ), .B1(_06609_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07378_ ) );
AOI22_X1 _22393_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06321_ ), .B1(_06360_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07379_ ) );
AOI21_X1 _22394_ ( .A(_06565_ ), .B1(_07378_ ), .B2(_07379_ ), .ZN(_07380_ ) );
OAI21_X1 _22395_ ( .A(_10261_ ), .B1(_07377_ ), .B2(_07380_ ), .ZN(_07381_ ) );
AOI22_X1 _22396_ ( .A1(_06580_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06325_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07382_ ) );
OAI211_X1 _22397_ ( .A(_06331_ ), .B(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06587_ ), .C2(_06588_ ), .ZN(_07383_ ) );
NAND3_X1 _22398_ ( .A1(_06925_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06249_ ), .ZN(_07384_ ) );
NAND4_X1 _22399_ ( .A1(_07382_ ), .A2(_06556_ ), .A3(_07383_ ), .A4(_07384_ ), .ZN(_07385_ ) );
AOI22_X1 _22400_ ( .A1(_06574_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06757_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07386_ ) );
AOI22_X1 _22401_ ( .A1(_06580_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06340_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07387_ ) );
NAND3_X1 _22402_ ( .A1(_07386_ ), .A2(_07387_ ), .A3(_06582_ ), .ZN(_07388_ ) );
NAND3_X1 _22403_ ( .A1(_06555_ ), .A2(_07385_ ), .A3(_07388_ ), .ZN(_07389_ ) );
NAND3_X1 _22404_ ( .A1(_07381_ ), .A2(_11056_ ), .A3(_07389_ ), .ZN(_07390_ ) );
NAND3_X1 _22405_ ( .A1(_07374_ ), .A2(_09805_ ), .A3(_07390_ ), .ZN(_07391_ ) );
NAND3_X1 _22406_ ( .A1(_07353_ ), .A2(_07391_ ), .A3(_09491_ ), .ZN(_07392_ ) );
AND3_X1 _22407_ ( .A1(_06557_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06678_ ), .ZN(_07393_ ) );
AOI221_X4 _22408_ ( .A(_07393_ ), .B1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06559_ ), .C1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06232_ ), .ZN(_07394_ ) );
NAND3_X1 _22409_ ( .A1(_06235_ ), .A2(_06562_ ), .A3(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07395_ ) );
NAND3_X1 _22410_ ( .A1(_07394_ ), .A2(_06576_ ), .A3(_07395_ ), .ZN(_07396_ ) );
AND3_X1 _22411_ ( .A1(_06239_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06256_ ), .ZN(_07397_ ) );
AOI221_X4 _22412_ ( .A(_07397_ ), .B1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06242_ ), .C1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C2(_06383_ ), .ZN(_07398_ ) );
NAND3_X1 _22413_ ( .A1(_06246_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06249_ ), .ZN(_07399_ ) );
NAND3_X1 _22414_ ( .A1(_07398_ ), .A2(_06245_ ), .A3(_07399_ ), .ZN(_07400_ ) );
AOI21_X1 _22415_ ( .A(_06463_ ), .B1(_07396_ ), .B2(_07400_ ), .ZN(_07401_ ) );
OAI211_X1 _22416_ ( .A(_06187_ ), .B(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(_05868_ ), .C2(_05869_ ), .ZN(_07402_ ) );
INV_X1 _22417_ ( .A(_07402_ ), .ZN(_07403_ ) );
AOI221_X4 _22418_ ( .A(_07403_ ), .B1(_06923_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .C2(_09626_ ), .ZN(_07404_ ) );
NAND3_X1 _22419_ ( .A1(_06473_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06333_ ), .ZN(_07405_ ) );
AOI21_X1 _22420_ ( .A(_06390_ ), .B1(_07404_ ), .B2(_07405_ ), .ZN(_07406_ ) );
AOI22_X1 _22421_ ( .A1(_06286_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06179_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07407_ ) );
AOI22_X1 _22422_ ( .A1(_06527_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06506_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07408_ ) );
AOI21_X1 _22423_ ( .A(_09084_ ), .B1(_07407_ ), .B2(_07408_ ), .ZN(_07409_ ) );
NOR3_X1 _22424_ ( .A1(_07406_ ), .A2(_06500_ ), .A3(_07409_ ), .ZN(_07410_ ) );
NOR3_X1 _22425_ ( .A1(_07401_ ), .A2(_07410_ ), .A3(_11196_ ), .ZN(_07411_ ) );
AOI22_X1 _22426_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06637_ ), .B1(_06366_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07412_ ) );
AOI22_X1 _22427_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06369_ ), .B1(_06370_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07413_ ) );
AOI21_X1 _22428_ ( .A(_06144_ ), .B1(_07412_ ), .B2(_07413_ ), .ZN(_07414_ ) );
AOI22_X1 _22429_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_09746_ ), .B1(_06429_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07415_ ) );
AOI22_X1 _22430_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06872_ ), .B1(_06864_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07416_ ) );
AOI21_X1 _22431_ ( .A(_06636_ ), .B1(_07415_ ), .B2(_07416_ ), .ZN(_07417_ ) );
OAI21_X1 _22432_ ( .A(_06645_ ), .B1(_07414_ ), .B2(_07417_ ), .ZN(_07418_ ) );
AOI22_X1 _22433_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06365_ ), .B1(_06263_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07419_ ) );
AOI22_X1 _22434_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06594_ ), .B1(_06370_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07420_ ) );
NAND3_X1 _22435_ ( .A1(_07419_ ), .A2(_06368_ ), .A3(_07420_ ), .ZN(_07421_ ) );
AOI22_X1 _22436_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06637_ ), .B1(_06366_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07422_ ) );
AOI22_X1 _22437_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06794_ ), .B1(_06702_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07423_ ) );
NAND3_X1 _22438_ ( .A1(_07422_ ), .A2(_06362_ ), .A3(_07423_ ), .ZN(_07424_ ) );
NAND3_X1 _22439_ ( .A1(_09056_ ), .A2(_07421_ ), .A3(_07424_ ), .ZN(_07425_ ) );
AOI21_X1 _22440_ ( .A(_09594_ ), .B1(_07418_ ), .B2(_07425_ ), .ZN(_07426_ ) );
OAI21_X1 _22441_ ( .A(_09489_ ), .B1(_07411_ ), .B2(_07426_ ), .ZN(_07427_ ) );
NAND3_X1 _22442_ ( .A1(_06671_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06399_ ), .ZN(_07428_ ) );
INV_X1 _22443_ ( .A(_07428_ ), .ZN(_07429_ ) );
AOI221_X4 _22444_ ( .A(_07429_ ), .B1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06430_ ), .C1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06326_ ), .ZN(_07430_ ) );
NAND3_X1 _22445_ ( .A1(_06561_ ), .A2(_06562_ ), .A3(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07431_ ) );
AOI21_X1 _22446_ ( .A(_06308_ ), .B1(_07430_ ), .B2(_07431_ ), .ZN(_07432_ ) );
NAND3_X1 _22447_ ( .A1(_06145_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06296_ ), .ZN(_07433_ ) );
INV_X1 _22448_ ( .A(_07433_ ), .ZN(_07434_ ) );
AOI221_X4 _22449_ ( .A(_07434_ ), .B1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06149_ ), .C1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06424_ ), .ZN(_07435_ ) );
NAND3_X1 _22450_ ( .A1(_06619_ ), .A2(_06569_ ), .A3(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07436_ ) );
AOI21_X1 _22451_ ( .A(_06209_ ), .B1(_07435_ ), .B2(_07436_ ), .ZN(_07437_ ) );
OAI21_X1 _22452_ ( .A(_06573_ ), .B1(_07432_ ), .B2(_07437_ ), .ZN(_07438_ ) );
AOI22_X1 _22453_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06305_ ), .B1(_06469_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07439_ ) );
AOI22_X1 _22454_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06757_ ), .B1(_06340_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07440_ ) );
NAND3_X1 _22455_ ( .A1(_07439_ ), .A2(_06582_ ), .A3(_07440_ ), .ZN(_07441_ ) );
AOI22_X1 _22456_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06305_ ), .B1(_06469_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07442_ ) );
AOI22_X1 _22457_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06757_ ), .B1(_06306_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07443_ ) );
NAND3_X1 _22458_ ( .A1(_07442_ ), .A2(_06576_ ), .A3(_07443_ ), .ZN(_07444_ ) );
NAND3_X1 _22459_ ( .A1(_06555_ ), .A2(_07441_ ), .A3(_07444_ ), .ZN(_07445_ ) );
NAND3_X1 _22460_ ( .A1(_07438_ ), .A2(_10053_ ), .A3(_07445_ ), .ZN(_07446_ ) );
AOI22_X1 _22461_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06205_ ), .B1(_06217_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07447_ ) );
AOI22_X1 _22462_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06220_ ), .B1(_06213_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07448_ ) );
NAND3_X1 _22463_ ( .A1(_07447_ ), .A2(_06209_ ), .A3(_07448_ ), .ZN(_07449_ ) );
AOI22_X1 _22464_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06216_ ), .B1(_06649_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07450_ ) );
AOI22_X1 _22465_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06347_ ), .B1(_06640_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07451_ ) );
NAND3_X1 _22466_ ( .A1(_07450_ ), .A2(_06964_ ), .A3(_07451_ ), .ZN(_07452_ ) );
NAND3_X1 _22467_ ( .A1(_06254_ ), .A2(_07449_ ), .A3(_07452_ ), .ZN(_07453_ ) );
AOI22_X1 _22468_ ( .A1(_06266_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06150_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07454_ ) );
OAI211_X1 _22469_ ( .A(_06436_ ), .B(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06352_ ), .C2(_06355_ ), .ZN(_07455_ ) );
NAND3_X1 _22470_ ( .A1(_06397_ ), .A2(_06598_ ), .A3(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07456_ ) );
AND3_X1 _22471_ ( .A1(_07454_ ), .A2(_07455_ ), .A3(_07456_ ), .ZN(_07457_ ) );
AOI22_X1 _22472_ ( .A1(_06266_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06150_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07458_ ) );
NAND3_X1 _22473_ ( .A1(_07362_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06797_ ), .ZN(_07459_ ) );
NAND3_X1 _22474_ ( .A1(_06397_ ), .A2(_06598_ ), .A3(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07460_ ) );
AND3_X1 _22475_ ( .A1(_07458_ ), .A2(_07459_ ), .A3(_07460_ ), .ZN(_07461_ ) );
MUX2_X1 _22476_ ( .A(_07457_ ), .B(_07461_ ), .S(_06433_ ), .Z(_07462_ ) );
OAI211_X1 _22477_ ( .A(_11196_ ), .B(_07453_ ), .C1(_07462_ ), .C2(_10261_ ), .ZN(_07463_ ) );
NAND3_X1 _22478_ ( .A1(_07446_ ), .A2(_06143_ ), .A3(_07463_ ), .ZN(_07464_ ) );
NAND3_X1 _22479_ ( .A1(_07427_ ), .A2(_02457_ ), .A3(_07464_ ), .ZN(_07465_ ) );
NAND3_X1 _22480_ ( .A1(_07392_ ), .A2(_09035_ ), .A3(_07465_ ), .ZN(_07466_ ) );
AND3_X1 _22481_ ( .A1(_06228_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06229_ ), .ZN(_07467_ ) );
AOI221_X4 _22482_ ( .A(_07467_ ), .B1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06231_ ), .C1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06285_ ), .ZN(_07468_ ) );
NAND3_X1 _22483_ ( .A1(_06568_ ), .A2(_06569_ ), .A3(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07469_ ) );
NAND3_X1 _22484_ ( .A1(_07468_ ), .A2(_06611_ ), .A3(_07469_ ), .ZN(_07470_ ) );
MUX2_X1 _22485_ ( .A(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .S(_06722_ ), .Z(_07471_ ) );
MUX2_X1 _22486_ ( .A(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .S(_06722_ ), .Z(_07472_ ) );
MUX2_X1 _22487_ ( .A(_07471_ ), .B(_07472_ ), .S(_06441_ ), .Z(_07473_ ) );
OAI211_X1 _22488_ ( .A(_07470_ ), .B(_09056_ ), .C1(_06721_ ), .C2(_07473_ ), .ZN(_07474_ ) );
AND3_X1 _22489_ ( .A1(_06439_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06296_ ), .ZN(_07475_ ) );
AOI221_X4 _22490_ ( .A(_07475_ ), .B1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06163_ ), .C1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .C2(_06206_ ), .ZN(_07476_ ) );
NAND3_X1 _22491_ ( .A1(_06718_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06675_ ), .ZN(_07477_ ) );
NAND3_X1 _22492_ ( .A1(_07476_ ), .A2(_06576_ ), .A3(_07477_ ), .ZN(_07478_ ) );
AND3_X1 _22493_ ( .A1(_06557_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06678_ ), .ZN(_07479_ ) );
AOI221_X4 _22494_ ( .A(_07479_ ), .B1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06559_ ), .C1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06266_ ), .ZN(_07480_ ) );
NAND3_X1 _22495_ ( .A1(_06561_ ), .A2(_06562_ ), .A3(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07481_ ) );
NAND3_X1 _22496_ ( .A1(_07480_ ), .A2(_06582_ ), .A3(_07481_ ), .ZN(_07482_ ) );
NAND3_X1 _22497_ ( .A1(_07478_ ), .A2(_07482_ ), .A3(_06315_ ), .ZN(_07483_ ) );
NAND3_X1 _22498_ ( .A1(_07474_ ), .A2(_07483_ ), .A3(_10053_ ), .ZN(_07484_ ) );
MUX2_X1 _22499_ ( .A(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .S(_06247_ ), .Z(_07485_ ) );
MUX2_X1 _22500_ ( .A(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .S(_06247_ ), .Z(_07486_ ) );
MUX2_X1 _22501_ ( .A(_07485_ ), .B(_07486_ ), .S(_10431_ ), .Z(_07487_ ) );
OAI21_X1 _22502_ ( .A(_09550_ ), .B1(_07487_ ), .B2(_06320_ ), .ZN(_07488_ ) );
AOI21_X1 _22503_ ( .A(_09119_ ), .B1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B2(_06384_ ), .ZN(_07489_ ) );
NAND3_X1 _22504_ ( .A1(_06441_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06408_ ), .ZN(_07490_ ) );
AOI22_X1 _22505_ ( .A1(_06177_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06506_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07491_ ) );
AND3_X1 _22506_ ( .A1(_07489_ ), .A2(_07490_ ), .A3(_07491_ ), .ZN(_07492_ ) );
AND3_X1 _22507_ ( .A1(_10430_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06392_ ), .ZN(_07493_ ) );
NAND3_X1 _22508_ ( .A1(_06434_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06543_ ), .ZN(_07494_ ) );
OAI211_X1 _22509_ ( .A(_06722_ ), .B(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06351_ ), .C2(_06354_ ), .ZN(_07495_ ) );
NAND2_X1 _22510_ ( .A1(_07494_ ), .A2(_07495_ ), .ZN(_07496_ ) );
AND3_X1 _22511_ ( .A1(_09069_ ), .A2(_09093_ ), .A3(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07497_ ) );
NOR3_X1 _22512_ ( .A1(_07493_ ), .A2(_07496_ ), .A3(_07497_ ), .ZN(_07498_ ) );
AND3_X1 _22513_ ( .A1(_06440_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06436_ ), .ZN(_07499_ ) );
OAI211_X1 _22514_ ( .A(_09093_ ), .B(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06351_ ), .C2(_06354_ ), .ZN(_07500_ ) );
NAND3_X1 _22515_ ( .A1(_09069_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06543_ ), .ZN(_07501_ ) );
NAND2_X1 _22516_ ( .A1(_07500_ ), .A2(_07501_ ), .ZN(_07502_ ) );
AND3_X1 _22517_ ( .A1(_09069_ ), .A2(_09093_ ), .A3(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07503_ ) );
NOR3_X1 _22518_ ( .A1(_07499_ ), .A2(_07502_ ), .A3(_07503_ ), .ZN(_07504_ ) );
MUX2_X1 _22519_ ( .A(_07498_ ), .B(_07504_ ), .S(_06495_ ), .Z(_07505_ ) );
OAI221_X1 _22520_ ( .A(_09665_ ), .B1(_07488_ ), .B2(_07492_ ), .C1(_07505_ ), .C2(_09744_ ), .ZN(_07506_ ) );
NAND3_X1 _22521_ ( .A1(_07484_ ), .A2(_06143_ ), .A3(_07506_ ), .ZN(_07507_ ) );
AND3_X1 _22522_ ( .A1(_06159_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_05809_ ), .ZN(_07508_ ) );
AOI221_X4 _22523_ ( .A(_07508_ ), .B1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06178_ ), .C1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06259_ ), .ZN(_07509_ ) );
NAND3_X1 _22524_ ( .A1(_06483_ ), .A2(_06599_ ), .A3(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07510_ ) );
NAND3_X1 _22525_ ( .A1(_07509_ ), .A2(_06514_ ), .A3(_07510_ ), .ZN(_07511_ ) );
MUX2_X1 _22526_ ( .A(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .S(_06247_ ), .Z(_07512_ ) );
MUX2_X1 _22527_ ( .A(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .S(_06199_ ), .Z(_07513_ ) );
MUX2_X1 _22528_ ( .A(_07512_ ), .B(_07513_ ), .S(_10431_ ), .Z(_07514_ ) );
OAI211_X1 _22529_ ( .A(_07511_ ), .B(_06500_ ), .C1(_09085_ ), .C2(_07514_ ), .ZN(_07515_ ) );
AOI22_X1 _22530_ ( .A1(_06343_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06422_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07516_ ) );
OAI211_X1 _22531_ ( .A(_06978_ ), .B(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06394_ ), .C2(_06395_ ), .ZN(_07517_ ) );
NAND3_X1 _22532_ ( .A1(_06398_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06401_ ), .ZN(_07518_ ) );
NAND4_X1 _22533_ ( .A1(_07516_ ), .A2(_06636_ ), .A3(_07517_ ), .A4(_07518_ ), .ZN(_07519_ ) );
AOI22_X1 _22534_ ( .A1(_06637_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06638_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07520_ ) );
AOI22_X1 _22535_ ( .A1(_06343_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06640_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07521_ ) );
NAND3_X1 _22536_ ( .A1(_07520_ ), .A2(_07521_ ), .A3(_06144_ ), .ZN(_07522_ ) );
NAND3_X1 _22537_ ( .A1(_06254_ ), .A2(_07519_ ), .A3(_07522_ ), .ZN(_07523_ ) );
AOI21_X1 _22538_ ( .A(_06413_ ), .B1(_07515_ ), .B2(_07523_ ), .ZN(_07524_ ) );
AOI22_X1 _22539_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06267_ ), .B1(_09795_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07525_ ) );
AOI22_X1 _22540_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06914_ ), .B1(_06915_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07526_ ) );
AOI21_X1 _22541_ ( .A(_07031_ ), .B1(_07525_ ), .B2(_07526_ ), .ZN(_07527_ ) );
AOI22_X1 _22542_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06286_ ), .B1(_06181_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07528_ ) );
AOI22_X1 _22543_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06264_ ), .B1(_06289_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07529_ ) );
AOI21_X1 _22544_ ( .A(_06284_ ), .B1(_07528_ ), .B2(_07529_ ), .ZN(_07530_ ) );
OAI21_X1 _22545_ ( .A(_06414_ ), .B1(_07527_ ), .B2(_07530_ ), .ZN(_07531_ ) );
AOI22_X1 _22546_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06286_ ), .B1(_06527_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07532_ ) );
AOI22_X1 _22547_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06264_ ), .B1(_06445_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07533_ ) );
AOI21_X1 _22548_ ( .A(_06495_ ), .B1(_07532_ ), .B2(_07533_ ), .ZN(_07534_ ) );
AOI22_X1 _22549_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06177_ ), .B1(_06504_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07535_ ) );
AOI22_X1 _22550_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06431_ ), .B1(_06506_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07536_ ) );
AOI21_X1 _22551_ ( .A(_06284_ ), .B1(_07535_ ), .B2(_07536_ ), .ZN(_07537_ ) );
OAI21_X1 _22552_ ( .A(_06500_ ), .B1(_07534_ ), .B2(_07537_ ), .ZN(_07538_ ) );
AOI21_X1 _22553_ ( .A(_10252_ ), .B1(_07531_ ), .B2(_07538_ ), .ZN(_07539_ ) );
OAI21_X1 _22554_ ( .A(_06227_ ), .B1(_07524_ ), .B2(_07539_ ), .ZN(_07540_ ) );
AOI21_X1 _22555_ ( .A(_09020_ ), .B1(_07507_ ), .B2(_07540_ ), .ZN(_07541_ ) );
AND3_X1 _22556_ ( .A1(_06557_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06391_ ), .ZN(_07542_ ) );
AOI221_X4 _22557_ ( .A(_07542_ ), .B1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06430_ ), .C1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C2(_06206_ ), .ZN(_07543_ ) );
NAND3_X1 _22558_ ( .A1(_06561_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06675_ ), .ZN(_07544_ ) );
NAND3_X1 _22559_ ( .A1(_07543_ ), .A2(_06300_ ), .A3(_07544_ ), .ZN(_07545_ ) );
AOI22_X1 _22560_ ( .A1(_06346_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06327_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07546_ ) );
NAND3_X1 _22561_ ( .A1(_06725_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06783_ ), .ZN(_07547_ ) );
NAND3_X1 _22562_ ( .A1(_06330_ ), .A2(_06331_ ), .A3(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07548_ ) );
NAND4_X1 _22563_ ( .A1(_07546_ ), .A2(_06329_ ), .A3(_07547_ ), .A4(_07548_ ), .ZN(_07549_ ) );
NAND3_X1 _22564_ ( .A1(_07545_ ), .A2(_10050_ ), .A3(_07549_ ), .ZN(_07550_ ) );
AOI22_X1 _22565_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06379_ ), .B1(_06380_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07551_ ) );
NAND3_X1 _22566_ ( .A1(_06473_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06333_ ), .ZN(_07552_ ) );
NAND3_X1 _22567_ ( .A1(_06483_ ), .A2(_06515_ ), .A3(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07553_ ) );
NAND4_X1 _22568_ ( .A1(_07551_ ), .A2(_06192_ ), .A3(_07552_ ), .A4(_07553_ ), .ZN(_07554_ ) );
AOI22_X1 _22569_ ( .A1(_06476_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06477_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07555_ ) );
NAND3_X1 _22570_ ( .A1(_06483_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06333_ ), .ZN(_07556_ ) );
OAI211_X1 _22571_ ( .A(_06939_ ), .B(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06480_ ), .C2(_06481_ ), .ZN(_07557_ ) );
NAND4_X1 _22572_ ( .A1(_07555_ ), .A2(_06700_ ), .A3(_07556_ ), .A4(_07557_ ), .ZN(_07558_ ) );
NAND3_X1 _22573_ ( .A1(_06645_ ), .A2(_07554_ ), .A3(_07558_ ), .ZN(_07559_ ) );
NAND3_X1 _22574_ ( .A1(_07550_ ), .A2(_09487_ ), .A3(_07559_ ), .ZN(_07560_ ) );
AOI22_X1 _22575_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06857_ ), .B1(_06343_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07561_ ) );
AOI22_X1 _22576_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06379_ ), .B1(_06380_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07562_ ) );
NAND3_X1 _22577_ ( .A1(_07561_ ), .A2(_06596_ ), .A3(_07562_ ), .ZN(_07563_ ) );
AOI22_X1 _22578_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06697_ ), .B1(_06360_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07564_ ) );
AOI22_X1 _22579_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06216_ ), .B1(_06649_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07565_ ) );
NAND3_X1 _22580_ ( .A1(_07564_ ), .A2(_06362_ ), .A3(_07565_ ), .ZN(_07566_ ) );
NAND3_X1 _22581_ ( .A1(_06645_ ), .A2(_07563_ ), .A3(_07566_ ), .ZN(_07567_ ) );
AOI22_X1 _22582_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06205_ ), .B1(_06217_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07568_ ) );
AOI22_X1 _22583_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06211_ ), .B1(_06213_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07569_ ) );
NAND3_X1 _22584_ ( .A1(_07568_ ), .A2(_06209_ ), .A3(_07569_ ), .ZN(_07570_ ) );
AOI22_X1 _22585_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06872_ ), .B1(_06640_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07571_ ) );
NAND3_X1 _22586_ ( .A1(_06492_ ), .A2(_06167_ ), .A3(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07572_ ) );
NAND3_X1 _22587_ ( .A1(_06398_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06931_ ), .ZN(_07573_ ) );
NAND4_X1 _22588_ ( .A1(_07571_ ), .A2(_06255_ ), .A3(_07572_ ), .A4(_07573_ ), .ZN(_07574_ ) );
NAND3_X1 _22589_ ( .A1(_06684_ ), .A2(_07570_ ), .A3(_07574_ ), .ZN(_07575_ ) );
NAND3_X1 _22590_ ( .A1(_07567_ ), .A2(_11196_ ), .A3(_07575_ ), .ZN(_07576_ ) );
NAND3_X1 _22591_ ( .A1(_07560_ ), .A2(_06338_ ), .A3(_07576_ ), .ZN(_07577_ ) );
AOI22_X1 _22592_ ( .A1(_06342_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06872_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07578_ ) );
NAND3_X1 _22593_ ( .A1(_06193_ ), .A2(_06194_ ), .A3(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07579_ ) );
NAND3_X1 _22594_ ( .A1(_06725_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06599_ ), .ZN(_07580_ ) );
NAND4_X1 _22595_ ( .A1(_07578_ ), .A2(_06964_ ), .A3(_07579_ ), .A4(_07580_ ), .ZN(_07581_ ) );
AOI22_X1 _22596_ ( .A1(_06365_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06380_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07582_ ) );
NAND3_X1 _22597_ ( .A1(_06473_ ), .A2(_06515_ ), .A3(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07583_ ) );
NAND3_X1 _22598_ ( .A1(_06725_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06484_ ), .ZN(_07584_ ) );
NAND4_X1 _22599_ ( .A1(_07582_ ), .A2(_06479_ ), .A3(_07583_ ), .A4(_07584_ ), .ZN(_07585_ ) );
NAND3_X1 _22600_ ( .A1(_06890_ ), .A2(_07581_ ), .A3(_07585_ ), .ZN(_07586_ ) );
AOI22_X1 _22601_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06325_ ), .B1(_06622_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07587_ ) );
AOI22_X1 _22602_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_09746_ ), .B1(_06540_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07588_ ) );
NAND3_X1 _22603_ ( .A1(_07587_ ), .A2(_06209_ ), .A3(_07588_ ), .ZN(_07589_ ) );
AOI22_X1 _22604_ ( .A1(_06836_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_09484_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07590_ ) );
NAND3_X1 _22605_ ( .A1(_06492_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06798_ ), .ZN(_07591_ ) );
OAI211_X1 _22606_ ( .A(_06978_ ), .B(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06394_ ), .C2(_06395_ ), .ZN(_07592_ ) );
NAND4_X1 _22607_ ( .A1(_07590_ ), .A2(_06255_ ), .A3(_07591_ ), .A4(_07592_ ), .ZN(_07593_ ) );
NAND3_X1 _22608_ ( .A1(_06252_ ), .A2(_07589_ ), .A3(_07593_ ), .ZN(_07594_ ) );
NAND3_X1 _22609_ ( .A1(_07586_ ), .A2(_09594_ ), .A3(_07594_ ), .ZN(_07595_ ) );
AOI22_X1 _22610_ ( .A1(_06318_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06638_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07596_ ) );
OAI211_X1 _22611_ ( .A(_06939_ ), .B(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06480_ ), .C2(_06481_ ), .ZN(_07597_ ) );
NAND3_X1 _22612_ ( .A1(_06166_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06798_ ), .ZN(_07598_ ) );
NAND4_X1 _22613_ ( .A1(_07596_ ), .A2(_06700_ ), .A3(_07597_ ), .A4(_07598_ ), .ZN(_07599_ ) );
AOI22_X1 _22614_ ( .A1(_06857_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06872_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07600_ ) );
AOI22_X1 _22615_ ( .A1(_06476_ ), .A2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06702_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07601_ ) );
NAND3_X1 _22616_ ( .A1(_07600_ ), .A2(_07601_ ), .A3(_06219_ ), .ZN(_07602_ ) );
NAND3_X1 _22617_ ( .A1(_06204_ ), .A2(_07599_ ), .A3(_07602_ ), .ZN(_07603_ ) );
AOI22_X1 _22618_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06794_ ), .B1(_06702_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07604_ ) );
AOI22_X1 _22619_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_07061_ ), .B1(_07062_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07605_ ) );
NAND3_X1 _22620_ ( .A1(_07604_ ), .A2(_06192_ ), .A3(_07605_ ), .ZN(_07606_ ) );
AOI22_X1 _22621_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_09746_ ), .B1(_06540_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07607_ ) );
AOI22_X1 _22622_ ( .A1(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06470_ ), .B1(_06864_ ), .B2(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07608_ ) );
NAND3_X1 _22623_ ( .A1(_07607_ ), .A2(_06700_ ), .A3(_07608_ ), .ZN(_07609_ ) );
NAND3_X1 _22624_ ( .A1(_06684_ ), .A2(_07606_ ), .A3(_07609_ ), .ZN(_07610_ ) );
NAND3_X1 _22625_ ( .A1(_07603_ ), .A2(_11196_ ), .A3(_07610_ ), .ZN(_07611_ ) );
NAND3_X1 _22626_ ( .A1(_07595_ ), .A2(_07611_ ), .A3(_10009_ ), .ZN(_07612_ ) );
AOI21_X1 _22627_ ( .A(_09018_ ), .B1(_07577_ ), .B2(_07612_ ), .ZN(_07613_ ) );
OAI21_X1 _22628_ ( .A(_09138_ ), .B1(_07541_ ), .B2(_07613_ ), .ZN(_07614_ ) );
AND3_X1 _22629_ ( .A1(_07466_ ), .A2(_07614_ ), .A3(_05734_ ), .ZN(\load_data_out[3] ) );
INV_X1 _22630_ ( .A(\load_data_out[3] ), .ZN(_07615_ ) );
OAI21_X1 _22631_ ( .A(_07615_ ), .B1(_10433_ ), .B2(_06130_ ), .ZN(_07616_ ) );
AOI21_X1 _22632_ ( .A(_07316_ ), .B1(_07616_ ), .B2(_06102_ ), .ZN(_07617_ ) );
NOR2_X1 _22633_ ( .A1(_07617_ ), .A2(_06137_ ), .ZN(_00026_ ) );
OAI22_X1 _22634_ ( .A1(_09096_ ), .A2(_05731_ ), .B1(\pc_out[2] ), .B2(_08928_ ), .ZN(_07618_ ) );
AND3_X1 _22635_ ( .A1(_06439_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06146_ ), .ZN(_07619_ ) );
AOI221_X4 _22636_ ( .A(_07619_ ), .B1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06716_ ), .C1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06266_ ), .ZN(_07620_ ) );
NAND3_X1 _22637_ ( .A1(_06718_ ), .A2(_06562_ ), .A3(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07621_ ) );
AOI21_X1 _22638_ ( .A(_06556_ ), .B1(_07620_ ), .B2(_07621_ ), .ZN(_07622_ ) );
AND3_X1 _22639_ ( .A1(_06228_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06256_ ), .ZN(_07623_ ) );
AOI221_X4 _22640_ ( .A(_07623_ ), .B1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06231_ ), .C1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06285_ ), .ZN(_07624_ ) );
NAND3_X1 _22641_ ( .A1(_06568_ ), .A2(_06236_ ), .A3(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07625_ ) );
AOI21_X1 _22642_ ( .A(_06565_ ), .B1(_07624_ ), .B2(_07625_ ), .ZN(_07626_ ) );
OAI21_X1 _22643_ ( .A(_09744_ ), .B1(_07622_ ), .B2(_07626_ ), .ZN(_07627_ ) );
AOI22_X1 _22644_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06574_ ), .B1(_06781_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07628_ ) );
AOI22_X1 _22645_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06339_ ), .B1(_09530_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07629_ ) );
NAND3_X1 _22646_ ( .A1(_07628_ ), .A2(_06300_ ), .A3(_07629_ ), .ZN(_07630_ ) );
AOI22_X1 _22647_ ( .A1(_06305_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06379_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07631_ ) );
NAND3_X1 _22648_ ( .A1(_06925_ ), .A2(_06811_ ), .A3(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07632_ ) );
OAI211_X1 _22649_ ( .A(_06515_ ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06587_ ), .C2(_06588_ ), .ZN(_07633_ ) );
NAND4_X1 _22650_ ( .A1(_07631_ ), .A2(_06308_ ), .A3(_07632_ ), .A4(_07633_ ), .ZN(_07634_ ) );
NAND3_X1 _22651_ ( .A1(_10261_ ), .A2(_07630_ ), .A3(_07634_ ), .ZN(_07635_ ) );
AOI21_X1 _22652_ ( .A(_06654_ ), .B1(_07627_ ), .B2(_07635_ ), .ZN(_07636_ ) );
AOI22_X1 _22653_ ( .A1(_06580_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06379_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07637_ ) );
OAI211_X1 _22654_ ( .A(_06515_ ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06587_ ), .C2(_06588_ ), .ZN(_07638_ ) );
NAND3_X1 _22655_ ( .A1(_06152_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06590_ ), .ZN(_07639_ ) );
NAND4_X1 _22656_ ( .A1(_07637_ ), .A2(_06308_ ), .A3(_07638_ ), .A4(_07639_ ), .ZN(_07640_ ) );
AOI22_X1 _22657_ ( .A1(_06580_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06697_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07641_ ) );
AOI22_X1 _22658_ ( .A1(_06305_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06340_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07642_ ) );
NAND3_X1 _22659_ ( .A1(_07641_ ), .A2(_07642_ ), .A3(_06582_ ), .ZN(_07643_ ) );
NAND3_X1 _22660_ ( .A1(_06573_ ), .A2(_07640_ ), .A3(_07643_ ), .ZN(_07644_ ) );
AOI22_X1 _22661_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06605_ ), .B1(_06318_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07645_ ) );
AOI22_X1 _22662_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06321_ ), .B1(_06360_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07646_ ) );
NAND3_X1 _22663_ ( .A1(_07645_ ), .A2(_06320_ ), .A3(_07646_ ), .ZN(_07647_ ) );
AOI22_X1 _22664_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06346_ ), .B1(_06609_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07648_ ) );
AOI22_X1 _22665_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06325_ ), .B1(_06327_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07649_ ) );
NAND3_X1 _22666_ ( .A1(_07648_ ), .A2(_06611_ ), .A3(_07649_ ), .ZN(_07650_ ) );
NAND3_X1 _22667_ ( .A1(_06303_ ), .A2(_07647_ ), .A3(_07650_ ), .ZN(_07651_ ) );
AOI21_X1 _22668_ ( .A(_09594_ ), .B1(_07644_ ), .B2(_07651_ ), .ZN(_07652_ ) );
OAI21_X1 _22669_ ( .A(_09489_ ), .B1(_07636_ ), .B2(_07652_ ), .ZN(_07653_ ) );
NAND3_X1 _22670_ ( .A1(_06671_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06399_ ), .ZN(_07654_ ) );
INV_X1 _22671_ ( .A(_07654_ ), .ZN(_07655_ ) );
AOI221_X4 _22672_ ( .A(_07655_ ), .B1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06163_ ), .C1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C2(_06206_ ), .ZN(_07656_ ) );
NAND3_X1 _22673_ ( .A1(_10432_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06675_ ), .ZN(_07657_ ) );
NAND3_X1 _22674_ ( .A1(_07656_ ), .A2(_06300_ ), .A3(_07657_ ), .ZN(_07658_ ) );
AOI22_X1 _22675_ ( .A1(_06305_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06340_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07659_ ) );
NAND3_X1 _22676_ ( .A1(_06246_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06249_ ), .ZN(_07660_ ) );
NAND3_X1 _22677_ ( .A1(_06309_ ), .A2(_06154_ ), .A3(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07661_ ) );
NAND4_X1 _22678_ ( .A1(_07659_ ), .A2(_06556_ ), .A3(_07660_ ), .A4(_07661_ ), .ZN(_07662_ ) );
NAND3_X1 _22679_ ( .A1(_07658_ ), .A2(_06555_ ), .A3(_07662_ ), .ZN(_07663_ ) );
AOI22_X1 _22680_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06857_ ), .B1(_06343_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07664_ ) );
AOI22_X1 _22681_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06325_ ), .B1(_06622_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07665_ ) );
AOI21_X1 _22682_ ( .A(_06964_ ), .B1(_07664_ ), .B2(_07665_ ), .ZN(_07666_ ) );
AOI22_X1 _22683_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06216_ ), .B1(_06217_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07667_ ) );
AOI22_X1 _22684_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06211_ ), .B1(_06213_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07668_ ) );
AOI21_X1 _22685_ ( .A(_06950_ ), .B1(_07667_ ), .B2(_07668_ ), .ZN(_07669_ ) );
OAI21_X1 _22686_ ( .A(_06890_ ), .B1(_07666_ ), .B2(_07669_ ), .ZN(_07670_ ) );
AOI21_X1 _22687_ ( .A(_09487_ ), .B1(_07663_ ), .B2(_07670_ ), .ZN(_07671_ ) );
AOI22_X1 _22688_ ( .A1(_06781_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06211_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07672_ ) );
NAND3_X1 _22689_ ( .A1(_06625_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06311_ ), .ZN(_07673_ ) );
OAI211_X1 _22690_ ( .A(_06167_ ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06600_ ), .C2(_06601_ ), .ZN(_07674_ ) );
NAND4_X1 _22691_ ( .A1(_07672_ ), .A2(_06565_ ), .A3(_07673_ ), .A4(_07674_ ), .ZN(_07675_ ) );
AOI22_X1 _22692_ ( .A1(_06305_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06379_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07676_ ) );
AOI22_X1 _22693_ ( .A1(_06593_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06322_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07677_ ) );
NAND3_X1 _22694_ ( .A1(_07676_ ), .A2(_07677_ ), .A3(_06556_ ), .ZN(_07678_ ) );
NAND3_X1 _22695_ ( .A1(_06573_ ), .A2(_07675_ ), .A3(_07678_ ), .ZN(_07679_ ) );
AOI22_X1 _22696_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06216_ ), .B1(_06217_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07680_ ) );
AOI22_X1 _22697_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06211_ ), .B1(_06213_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07681_ ) );
AOI21_X1 _22698_ ( .A(_06950_ ), .B1(_07680_ ), .B2(_07681_ ), .ZN(_07682_ ) );
AOI22_X1 _22699_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06382_ ), .B1(_06384_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07683_ ) );
AOI22_X1 _22700_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06477_ ), .B1(_06425_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07684_ ) );
AOI21_X1 _22701_ ( .A(_07031_ ), .B1(_07683_ ), .B2(_07684_ ), .ZN(_07685_ ) );
OAI21_X1 _22702_ ( .A(_06252_ ), .B1(_07682_ ), .B2(_07685_ ), .ZN(_07686_ ) );
AOI21_X1 _22703_ ( .A(_11196_ ), .B1(_07679_ ), .B2(_07686_ ), .ZN(_07687_ ) );
OAI21_X1 _22704_ ( .A(_09805_ ), .B1(_07671_ ), .B2(_07687_ ), .ZN(_07688_ ) );
NAND3_X1 _22705_ ( .A1(_07653_ ), .A2(_07688_ ), .A3(_02409_ ), .ZN(_07689_ ) );
AND3_X1 _22706_ ( .A1(_06456_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06160_ ), .ZN(_07690_ ) );
AOI221_X4 _22707_ ( .A(_07690_ ), .B1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06923_ ), .C1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06176_ ), .ZN(_07691_ ) );
NAND3_X1 _22708_ ( .A1(_06152_ ), .A2(_06154_ ), .A3(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07692_ ) );
NAND3_X1 _22709_ ( .A1(_07691_ ), .A2(_06362_ ), .A3(_07692_ ), .ZN(_07693_ ) );
MUX2_X1 _22710_ ( .A(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .S(_06464_ ), .Z(_07694_ ) );
MUX2_X1 _22711_ ( .A(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .S(_06464_ ), .Z(_07695_ ) );
MUX2_X1 _22712_ ( .A(_07694_ ), .B(_07695_ ), .S(_06448_ ), .Z(_07696_ ) );
OAI211_X1 _22713_ ( .A(_07693_ ), .B(_06254_ ), .C1(_06198_ ), .C2(_07696_ ), .ZN(_07697_ ) );
AND3_X1 _22714_ ( .A1(_07362_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06400_ ), .ZN(_07698_ ) );
OAI211_X1 _22715_ ( .A(_06392_ ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06351_ ), .C2(_06354_ ), .ZN(_07699_ ) );
NAND3_X1 _22716_ ( .A1(_06434_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06436_ ), .ZN(_07700_ ) );
NAND2_X1 _22717_ ( .A1(_07699_ ), .A2(_07700_ ), .ZN(_07701_ ) );
AND3_X1 _22718_ ( .A1(_06434_ ), .A2(_06392_ ), .A3(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07702_ ) );
NOR3_X1 _22719_ ( .A1(_07698_ ), .A2(_07701_ ), .A3(_07702_ ), .ZN(_07703_ ) );
AOI22_X1 _22720_ ( .A1(_06298_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06424_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07704_ ) );
NAND3_X1 _22721_ ( .A1(_07362_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06797_ ), .ZN(_07705_ ) );
NAND3_X1 _22722_ ( .A1(_06397_ ), .A2(_06153_ ), .A3(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07706_ ) );
AND3_X1 _22723_ ( .A1(_07704_ ), .A2(_07705_ ), .A3(_07706_ ), .ZN(_07707_ ) );
MUX2_X1 _22724_ ( .A(_07703_ ), .B(_07707_ ), .S(_06158_ ), .Z(_07708_ ) );
OAI211_X1 _22725_ ( .A(_07697_ ), .B(_11056_ ), .C1(_10529_ ), .C2(_07708_ ), .ZN(_07709_ ) );
AND3_X1 _22726_ ( .A1(_06439_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06146_ ), .ZN(_07710_ ) );
AOI221_X4 _22727_ ( .A(_07710_ ), .B1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06716_ ), .C1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06266_ ), .ZN(_07711_ ) );
NAND3_X1 _22728_ ( .A1(_06718_ ), .A2(_09095_ ), .A3(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07712_ ) );
AOI21_X1 _22729_ ( .A(_06556_ ), .B1(_07711_ ), .B2(_07712_ ), .ZN(_07713_ ) );
AND3_X1 _22730_ ( .A1(_06228_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06256_ ), .ZN(_07714_ ) );
AOI221_X4 _22731_ ( .A(_07714_ ), .B1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06231_ ), .C1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .C2(_06383_ ), .ZN(_07715_ ) );
NAND3_X1 _22732_ ( .A1(_06568_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06736_ ), .ZN(_07716_ ) );
AOI21_X1 _22733_ ( .A(_06565_ ), .B1(_07715_ ), .B2(_07716_ ), .ZN(_07717_ ) );
OAI21_X1 _22734_ ( .A(_10261_ ), .B1(_07713_ ), .B2(_07717_ ), .ZN(_07718_ ) );
AND3_X1 _22735_ ( .A1(_06456_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06240_ ), .ZN(_07719_ ) );
AOI221_X4 _22736_ ( .A(_07719_ ), .B1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06242_ ), .C1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06176_ ), .ZN(_07720_ ) );
NAND3_X1 _22737_ ( .A1(_06619_ ), .A2(_06811_ ), .A3(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07721_ ) );
NAND3_X1 _22738_ ( .A1(_07720_ ), .A2(_06556_ ), .A3(_07721_ ), .ZN(_07722_ ) );
MUX2_X1 _22739_ ( .A(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .S(_06464_ ), .Z(_07723_ ) );
MUX2_X1 _22740_ ( .A(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .S(_06464_ ), .Z(_07724_ ) );
MUX2_X1 _22741_ ( .A(_07723_ ), .B(_07724_ ), .S(_06448_ ), .Z(_07725_ ) );
OAI211_X1 _22742_ ( .A(_07722_ ), .B(_06252_ ), .C1(_06721_ ), .C2(_07725_ ), .ZN(_07726_ ) );
NAND3_X1 _22743_ ( .A1(_07718_ ), .A2(_09784_ ), .A3(_07726_ ), .ZN(_07727_ ) );
NAND3_X1 _22744_ ( .A1(_07709_ ), .A2(_07727_ ), .A3(_06143_ ), .ZN(_07728_ ) );
AND3_X1 _22745_ ( .A1(_06239_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06229_ ), .ZN(_07729_ ) );
AOI221_X4 _22746_ ( .A(_07729_ ), .B1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06231_ ), .C1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .C2(_06383_ ), .ZN(_07730_ ) );
NAND3_X1 _22747_ ( .A1(_10432_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06736_ ), .ZN(_07731_ ) );
NAND3_X1 _22748_ ( .A1(_07730_ ), .A2(_06234_ ), .A3(_07731_ ), .ZN(_07732_ ) );
MUX2_X1 _22749_ ( .A(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .S(_06722_ ), .Z(_07733_ ) );
MUX2_X1 _22750_ ( .A(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .S(_06722_ ), .Z(_07734_ ) );
MUX2_X1 _22751_ ( .A(_07733_ ), .B(_07734_ ), .S(_06441_ ), .Z(_07735_ ) );
OAI211_X1 _22752_ ( .A(_07732_ ), .B(_10050_ ), .C1(_06721_ ), .C2(_07735_ ), .ZN(_07736_ ) );
AOI22_X1 _22753_ ( .A1(_06580_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06594_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07737_ ) );
NAND3_X1 _22754_ ( .A1(_06309_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06590_ ), .ZN(_07738_ ) );
OAI211_X1 _22755_ ( .A(_06599_ ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06587_ ), .C2(_06588_ ), .ZN(_07739_ ) );
NAND4_X1 _22756_ ( .A1(_07737_ ), .A2(_06596_ ), .A3(_07738_ ), .A4(_07739_ ), .ZN(_07740_ ) );
AOI22_X1 _22757_ ( .A1(_06593_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06369_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07741_ ) );
NAND3_X1 _22758_ ( .A1(_06459_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06311_ ), .ZN(_07742_ ) );
OAI211_X1 _22759_ ( .A(_06599_ ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06600_ ), .C2(_06601_ ), .ZN(_07743_ ) );
NAND4_X1 _22760_ ( .A1(_07741_ ), .A2(_06362_ ), .A3(_07742_ ), .A4(_07743_ ), .ZN(_07744_ ) );
NAND3_X1 _22761_ ( .A1(_06573_ ), .A2(_07740_ ), .A3(_07744_ ), .ZN(_07745_ ) );
NAND3_X1 _22762_ ( .A1(_07736_ ), .A2(_10053_ ), .A3(_07745_ ), .ZN(_07746_ ) );
AOI22_X1 _22763_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06605_ ), .B1(_06609_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07747_ ) );
AOI22_X1 _22764_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06697_ ), .B1(_06327_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07748_ ) );
AOI21_X1 _22765_ ( .A(_06329_ ), .B1(_07747_ ), .B2(_07748_ ), .ZN(_07749_ ) );
AOI22_X1 _22766_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06637_ ), .B1(_06207_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07750_ ) );
AOI22_X1 _22767_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06794_ ), .B1(_06702_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07751_ ) );
AOI21_X1 _22768_ ( .A(_06700_ ), .B1(_07750_ ), .B2(_07751_ ), .ZN(_07752_ ) );
OAI21_X1 _22769_ ( .A(_06315_ ), .B1(_07749_ ), .B2(_07752_ ), .ZN(_07753_ ) );
AOI22_X1 _22770_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06365_ ), .B1(_06366_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07754_ ) );
AOI22_X1 _22771_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06594_ ), .B1(_06370_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07755_ ) );
AOI21_X1 _22772_ ( .A(_06144_ ), .B1(_07754_ ), .B2(_07755_ ), .ZN(_07756_ ) );
AOI22_X1 _22773_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_09746_ ), .B1(_06429_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07757_ ) );
AOI22_X1 _22774_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06872_ ), .B1(_06864_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07758_ ) );
AOI21_X1 _22775_ ( .A(_06636_ ), .B1(_07757_ ), .B2(_07758_ ), .ZN(_07759_ ) );
OAI21_X1 _22776_ ( .A(_09056_ ), .B1(_07756_ ), .B2(_07759_ ), .ZN(_07760_ ) );
NAND3_X1 _22777_ ( .A1(_07753_ ), .A2(_06654_ ), .A3(_07760_ ), .ZN(_07761_ ) );
NAND3_X1 _22778_ ( .A1(_07746_ ), .A2(_10744_ ), .A3(_07761_ ), .ZN(_07762_ ) );
NAND3_X1 _22779_ ( .A1(_07728_ ), .A2(_09604_ ), .A3(_07762_ ), .ZN(_07763_ ) );
NAND3_X1 _22780_ ( .A1(_07689_ ), .A2(_09035_ ), .A3(_07763_ ), .ZN(_07764_ ) );
AND3_X1 _22781_ ( .A1(_06557_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06391_ ), .ZN(_07765_ ) );
AOI221_X4 _22782_ ( .A(_07765_ ), .B1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06430_ ), .C1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C2(_06383_ ), .ZN(_07766_ ) );
NAND3_X1 _22783_ ( .A1(_06235_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06736_ ), .ZN(_07767_ ) );
NAND3_X1 _22784_ ( .A1(_07766_ ), .A2(_06582_ ), .A3(_07767_ ), .ZN(_07768_ ) );
AOI22_X1 _22785_ ( .A1(_06857_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06622_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07769_ ) );
NAND3_X1 _22786_ ( .A1(_06725_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06783_ ), .ZN(_07770_ ) );
NAND3_X1 _22787_ ( .A1(_06473_ ), .A2(_06515_ ), .A3(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07771_ ) );
NAND4_X1 _22788_ ( .A1(_07769_ ), .A2(_06964_ ), .A3(_07770_ ), .A4(_07771_ ), .ZN(_07772_ ) );
NAND3_X1 _22789_ ( .A1(_07768_ ), .A2(_09056_ ), .A3(_07772_ ), .ZN(_07773_ ) );
AOI22_X1 _22790_ ( .A1(_06476_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06477_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07774_ ) );
OAI211_X1 _22791_ ( .A(_06350_ ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06480_ ), .C2(_06481_ ), .ZN(_07775_ ) );
NAND3_X1 _22792_ ( .A1(_06166_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06484_ ), .ZN(_07776_ ) );
NAND4_X1 _22793_ ( .A1(_07774_ ), .A2(_06700_ ), .A3(_07775_ ), .A4(_07776_ ), .ZN(_07777_ ) );
AOI22_X1 _22794_ ( .A1(_06346_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06220_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07778_ ) );
AOI22_X1 _22795_ ( .A1(_06476_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06370_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07779_ ) );
NAND3_X1 _22796_ ( .A1(_07778_ ), .A2(_07779_ ), .A3(_06329_ ), .ZN(_07780_ ) );
NAND3_X1 _22797_ ( .A1(_06645_ ), .A2(_07777_ ), .A3(_07780_ ), .ZN(_07781_ ) );
AOI21_X1 _22798_ ( .A(_11196_ ), .B1(_07773_ ), .B2(_07781_ ), .ZN(_07782_ ) );
AOI22_X1 _22799_ ( .A1(_06343_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06422_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07783_ ) );
OAI211_X1 _22800_ ( .A(_06978_ ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06394_ ), .C2(_06395_ ), .ZN(_07784_ ) );
NAND3_X1 _22801_ ( .A1(_06398_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06401_ ), .ZN(_07785_ ) );
NAND4_X1 _22802_ ( .A1(_07783_ ), .A2(_06405_ ), .A3(_07784_ ), .A4(_07785_ ), .ZN(_07786_ ) );
AOI22_X1 _22803_ ( .A1(_06609_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06914_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07787_ ) );
AOI22_X1 _22804_ ( .A1(_06421_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06864_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07788_ ) );
NAND3_X1 _22805_ ( .A1(_07787_ ), .A2(_07788_ ), .A3(_06973_ ), .ZN(_07789_ ) );
NAND3_X1 _22806_ ( .A1(_06463_ ), .A2(_07786_ ), .A3(_07789_ ), .ZN(_07790_ ) );
AOI22_X1 _22807_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06347_ ), .B1(_06640_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07791_ ) );
AOI22_X1 _22808_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06444_ ), .B1(_06527_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07792_ ) );
NAND3_X1 _22809_ ( .A1(_07791_ ), .A2(_06929_ ), .A3(_07792_ ), .ZN(_07793_ ) );
AOI22_X1 _22810_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_07061_ ), .B1(_09795_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07794_ ) );
AOI22_X1 _22811_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06914_ ), .B1(_06268_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07795_ ) );
NAND3_X1 _22812_ ( .A1(_07794_ ), .A2(_06950_ ), .A3(_07795_ ), .ZN(_07796_ ) );
NAND3_X1 _22813_ ( .A1(_06388_ ), .A2(_07793_ ), .A3(_07796_ ), .ZN(_07797_ ) );
AOI21_X1 _22814_ ( .A(_10252_ ), .B1(_07790_ ), .B2(_07797_ ), .ZN(_07798_ ) );
NOR3_X1 _22815_ ( .A1(_07782_ ), .A2(_07798_ ), .A3(_10009_ ), .ZN(_07799_ ) );
AOI22_X1 _22816_ ( .A1(_06609_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06914_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07800_ ) );
OAI211_X1 _22817_ ( .A(_06939_ ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06480_ ), .C2(_06481_ ), .ZN(_07801_ ) );
NAND3_X1 _22818_ ( .A1(_06166_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06798_ ), .ZN(_07802_ ) );
NAND4_X1 _22819_ ( .A1(_07800_ ), .A2(_06973_ ), .A3(_07801_ ), .A4(_07802_ ), .ZN(_07803_ ) );
AOI22_X1 _22820_ ( .A1(_06342_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06872_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07804_ ) );
AOI22_X1 _22821_ ( .A1(_06476_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06274_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07805_ ) );
NAND3_X1 _22822_ ( .A1(_07804_ ), .A2(_07805_ ), .A3(_06964_ ), .ZN(_07806_ ) );
NAND3_X1 _22823_ ( .A1(_06204_ ), .A2(_07803_ ), .A3(_07806_ ), .ZN(_07807_ ) );
AOI22_X1 _22824_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06369_ ), .B1(_06702_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07808_ ) );
AOI22_X1 _22825_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_07061_ ), .B1(_07062_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07809_ ) );
NAND3_X1 _22826_ ( .A1(_07808_ ), .A2(_06192_ ), .A3(_07809_ ), .ZN(_07810_ ) );
AOI22_X1 _22827_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_09746_ ), .B1(_06429_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07811_ ) );
AOI22_X1 _22828_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06470_ ), .B1(_06864_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07812_ ) );
NAND3_X1 _22829_ ( .A1(_07811_ ), .A2(_06700_ ), .A3(_07812_ ), .ZN(_07813_ ) );
NAND3_X1 _22830_ ( .A1(_06684_ ), .A2(_07810_ ), .A3(_07813_ ), .ZN(_07814_ ) );
AOI21_X1 _22831_ ( .A(_06186_ ), .B1(_07807_ ), .B2(_07814_ ), .ZN(_07815_ ) );
AOI22_X1 _22832_ ( .A1(_06267_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06268_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07816_ ) );
NAND3_X1 _22833_ ( .A1(_06407_ ), .A2(_06978_ ), .A3(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07817_ ) );
NAND3_X1 _22834_ ( .A1(_06441_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06437_ ), .ZN(_07818_ ) );
NAND4_X1 _22835_ ( .A1(_07816_ ), .A2(_06158_ ), .A3(_07817_ ), .A4(_07818_ ), .ZN(_07819_ ) );
AOI22_X1 _22836_ ( .A1(_06444_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06445_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07820_ ) );
NAND3_X1 _22837_ ( .A1(_06435_ ), .A2(_06978_ ), .A3(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07821_ ) );
NAND3_X1 _22838_ ( .A1(_06448_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06437_ ), .ZN(_07822_ ) );
NAND4_X1 _22839_ ( .A1(_07820_ ), .A2(_06197_ ), .A3(_07821_ ), .A4(_07822_ ), .ZN(_07823_ ) );
NAND3_X1 _22840_ ( .A1(_09482_ ), .A2(_07819_ ), .A3(_07823_ ), .ZN(_07824_ ) );
AOI22_X1 _22841_ ( .A1(_06286_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06289_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07825_ ) );
OAI211_X1 _22842_ ( .A(_06544_ ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06417_ ), .C2(_06418_ ), .ZN(_07826_ ) );
NAND3_X1 _22843_ ( .A1(_09070_ ), .A2(_06393_ ), .A3(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07827_ ) );
NAND4_X1 _22844_ ( .A1(_07825_ ), .A2(_06284_ ), .A3(_07826_ ), .A4(_07827_ ), .ZN(_07828_ ) );
AOI22_X1 _22845_ ( .A1(_06267_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06288_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07829_ ) );
AOI22_X1 _22846_ ( .A1(_06384_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06289_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07830_ ) );
NAND3_X1 _22847_ ( .A1(_07829_ ), .A2(_07830_ ), .A3(_06197_ ), .ZN(_07831_ ) );
NAND3_X1 _22848_ ( .A1(_06500_ ), .A2(_07828_ ), .A3(_07831_ ), .ZN(_07832_ ) );
AOI21_X1 _22849_ ( .A(_06413_ ), .B1(_07824_ ), .B2(_07832_ ), .ZN(_07833_ ) );
NOR3_X1 _22850_ ( .A1(_07815_ ), .A2(_07833_ ), .A3(_08995_ ), .ZN(_07834_ ) );
OAI21_X1 _22851_ ( .A(_02457_ ), .B1(_07799_ ), .B2(_07834_ ), .ZN(_07835_ ) );
AND3_X1 _22852_ ( .A1(_06228_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06229_ ), .ZN(_07836_ ) );
AOI221_X4 _22853_ ( .A(_07836_ ), .B1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06231_ ), .C1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06232_ ), .ZN(_07837_ ) );
NAND3_X1 _22854_ ( .A1(_06235_ ), .A2(_06236_ ), .A3(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07838_ ) );
NAND3_X1 _22855_ ( .A1(_07837_ ), .A2(_06234_ ), .A3(_07838_ ), .ZN(_07839_ ) );
MUX2_X1 _22856_ ( .A(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .S(_06722_ ), .Z(_07840_ ) );
MUX2_X1 _22857_ ( .A(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .S(_06722_ ), .Z(_07841_ ) );
MUX2_X1 _22858_ ( .A(_07840_ ), .B(_07841_ ), .S(_06441_ ), .Z(_07842_ ) );
OAI211_X1 _22859_ ( .A(_07839_ ), .B(_09056_ ), .C1(_06721_ ), .C2(_07842_ ), .ZN(_07843_ ) );
AND3_X1 _22860_ ( .A1(_06439_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06296_ ), .ZN(_07844_ ) );
AOI221_X4 _22861_ ( .A(_07844_ ), .B1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06163_ ), .C1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06298_ ), .ZN(_07845_ ) );
NAND3_X1 _22862_ ( .A1(_06718_ ), .A2(_09095_ ), .A3(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07846_ ) );
NAND3_X1 _22863_ ( .A1(_07845_ ), .A2(_09085_ ), .A3(_07846_ ), .ZN(_07847_ ) );
AND3_X1 _22864_ ( .A1(_06439_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06146_ ), .ZN(_07848_ ) );
AOI221_X4 _22865_ ( .A(_07848_ ), .B1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06716_ ), .C1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C2(_06206_ ), .ZN(_07849_ ) );
NAND3_X1 _22866_ ( .A1(_06561_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06675_ ), .ZN(_07850_ ) );
NAND3_X1 _22867_ ( .A1(_07849_ ), .A2(_06300_ ), .A3(_07850_ ), .ZN(_07851_ ) );
NAND3_X1 _22868_ ( .A1(_07847_ ), .A2(_07851_ ), .A3(_06315_ ), .ZN(_07852_ ) );
NAND3_X1 _22869_ ( .A1(_07843_ ), .A2(_07852_ ), .A3(_10053_ ), .ZN(_07853_ ) );
MUX2_X1 _22870_ ( .A(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .S(_06247_ ), .Z(_07854_ ) );
MUX2_X1 _22871_ ( .A(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .S(_06247_ ), .Z(_07855_ ) );
MUX2_X1 _22872_ ( .A(_07854_ ), .B(_07855_ ), .S(_10431_ ), .Z(_07856_ ) );
OAI21_X1 _22873_ ( .A(_09550_ ), .B1(_07856_ ), .B2(_06320_ ), .ZN(_07857_ ) );
AOI21_X1 _22874_ ( .A(_09119_ ), .B1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B2(_06429_ ), .ZN(_07858_ ) );
NAND3_X1 _22875_ ( .A1(_06441_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06408_ ), .ZN(_07859_ ) );
AOI22_X1 _22876_ ( .A1(_06177_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06506_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07860_ ) );
AND3_X1 _22877_ ( .A1(_07858_ ), .A2(_07859_ ), .A3(_07860_ ), .ZN(_07861_ ) );
AND3_X1 _22878_ ( .A1(_06440_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06436_ ), .ZN(_07862_ ) );
OAI211_X1 _22879_ ( .A(_09093_ ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06351_ ), .C2(_06354_ ), .ZN(_07863_ ) );
NAND3_X1 _22880_ ( .A1(_09069_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06543_ ), .ZN(_07864_ ) );
NAND2_X1 _22881_ ( .A1(_07863_ ), .A2(_07864_ ), .ZN(_07865_ ) );
AND3_X1 _22882_ ( .A1(_09069_ ), .A2(_09093_ ), .A3(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07866_ ) );
NOR3_X1 _22883_ ( .A1(_07862_ ), .A2(_07865_ ), .A3(_07866_ ), .ZN(_07867_ ) );
AND3_X1 _22884_ ( .A1(_06440_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06436_ ), .ZN(_07868_ ) );
OAI211_X1 _22885_ ( .A(_06392_ ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06351_ ), .C2(_06354_ ), .ZN(_07869_ ) );
NAND3_X1 _22886_ ( .A1(_09069_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06543_ ), .ZN(_07870_ ) );
NAND2_X1 _22887_ ( .A1(_07869_ ), .A2(_07870_ ), .ZN(_07871_ ) );
AND3_X1 _22888_ ( .A1(_09069_ ), .A2(_06392_ ), .A3(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07872_ ) );
NOR3_X1 _22889_ ( .A1(_07868_ ), .A2(_07871_ ), .A3(_07872_ ), .ZN(_07873_ ) );
MUX2_X1 _22890_ ( .A(_07867_ ), .B(_07873_ ), .S(_06495_ ), .Z(_07874_ ) );
OAI221_X1 _22891_ ( .A(_09665_ ), .B1(_07857_ ), .B2(_07861_ ), .C1(_07874_ ), .C2(_09744_ ), .ZN(_07875_ ) );
NAND3_X1 _22892_ ( .A1(_07853_ ), .A2(_06143_ ), .A3(_07875_ ), .ZN(_07876_ ) );
AND3_X1 _22893_ ( .A1(_06159_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_05809_ ), .ZN(_07877_ ) );
AOI221_X4 _22894_ ( .A(_07877_ ), .B1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_09528_ ), .C1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .C2(_09626_ ), .ZN(_07878_ ) );
NAND3_X1 _22895_ ( .A1(_06725_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06333_ ), .ZN(_07879_ ) );
NAND3_X1 _22896_ ( .A1(_07878_ ), .A2(_06514_ ), .A3(_07879_ ), .ZN(_07880_ ) );
MUX2_X1 _22897_ ( .A(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .S(_06199_ ), .Z(_07881_ ) );
MUX2_X1 _22898_ ( .A(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .S(_06199_ ), .Z(_07882_ ) );
MUX2_X1 _22899_ ( .A(_07881_ ), .B(_07882_ ), .S(_10431_ ), .Z(_07883_ ) );
OAI211_X1 _22900_ ( .A(_07880_ ), .B(_06500_ ), .C1(_06198_ ), .C2(_07883_ ), .ZN(_07884_ ) );
AOI22_X1 _22901_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06216_ ), .B1(_06649_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07885_ ) );
AOI22_X1 _22902_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06220_ ), .B1(_06221_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07886_ ) );
NAND3_X1 _22903_ ( .A1(_07885_ ), .A2(_06479_ ), .A3(_07886_ ), .ZN(_07887_ ) );
AOI22_X1 _22904_ ( .A1(_06637_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06638_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_07888_ ) );
AOI22_X1 _22905_ ( .A1(_06836_ ), .A2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06221_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07889_ ) );
NAND3_X1 _22906_ ( .A1(_07888_ ), .A2(_07889_ ), .A3(_06144_ ), .ZN(_07890_ ) );
NAND3_X1 _22907_ ( .A1(_06254_ ), .A2(_07887_ ), .A3(_07890_ ), .ZN(_07891_ ) );
AOI21_X1 _22908_ ( .A(_06413_ ), .B1(_07884_ ), .B2(_07891_ ), .ZN(_07892_ ) );
AOI22_X1 _22909_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_07061_ ), .B1(_07062_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07893_ ) );
AOI22_X1 _22910_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06914_ ), .B1(_06915_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07894_ ) );
AOI21_X1 _22911_ ( .A(_07031_ ), .B1(_07893_ ), .B2(_07894_ ), .ZN(_07895_ ) );
AOI22_X1 _22912_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06286_ ), .B1(_06181_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07896_ ) );
AOI22_X1 _22913_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06264_ ), .B1(_06289_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07897_ ) );
AOI21_X1 _22914_ ( .A(_06284_ ), .B1(_07896_ ), .B2(_07897_ ), .ZN(_07898_ ) );
OAI21_X1 _22915_ ( .A(_06414_ ), .B1(_07895_ ), .B2(_07898_ ), .ZN(_07899_ ) );
AOI22_X1 _22916_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_07061_ ), .B1(_07062_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07900_ ) );
AOI22_X1 _22917_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06914_ ), .B1(_06915_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07901_ ) );
NAND3_X1 _22918_ ( .A1(_07900_ ), .A2(_06929_ ), .A3(_07901_ ), .ZN(_07902_ ) );
AOI22_X1 _22919_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06267_ ), .B1(_09795_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07903_ ) );
AOI22_X1 _22920_ ( .A1(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_09484_ ), .B1(_06268_ ), .B2(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07904_ ) );
NAND3_X1 _22921_ ( .A1(_07903_ ), .A2(_06950_ ), .A3(_07904_ ), .ZN(_07905_ ) );
NAND3_X1 _22922_ ( .A1(_09463_ ), .A2(_07902_ ), .A3(_07905_ ), .ZN(_07906_ ) );
AOI21_X1 _22923_ ( .A(_10252_ ), .B1(_07899_ ), .B2(_07906_ ), .ZN(_07907_ ) );
OAI21_X1 _22924_ ( .A(_06227_ ), .B1(_07892_ ), .B2(_07907_ ), .ZN(_07908_ ) );
NAND3_X1 _22925_ ( .A1(_07876_ ), .A2(_09604_ ), .A3(_07908_ ), .ZN(_07909_ ) );
NAND3_X1 _22926_ ( .A1(_07835_ ), .A2(_09138_ ), .A3(_07909_ ), .ZN(_07910_ ) );
AND3_X1 _22927_ ( .A1(_07764_ ), .A2(_06077_ ), .A3(_07910_ ), .ZN(\load_data_out[2] ) );
INV_X1 _22928_ ( .A(\load_data_out[2] ), .ZN(_07911_ ) );
OAI21_X1 _22929_ ( .A(_07911_ ), .B1(_09096_ ), .B2(_06130_ ), .ZN(_07912_ ) );
AOI21_X1 _22930_ ( .A(_07618_ ), .B1(_07912_ ), .B2(_06101_ ), .ZN(_07913_ ) );
NOR2_X1 _22931_ ( .A1(_07913_ ), .A2(_06137_ ), .ZN(_00027_ ) );
AND2_X1 _22932_ ( .A1(\alu_result_out[28] ), .A2(_06078_ ), .ZN(_07914_ ) );
OAI21_X1 _22933_ ( .A(_06065_ ), .B1(_06077_ ), .B2(_07914_ ), .ZN(_07915_ ) );
AOI22_X1 _22934_ ( .A1(\alu_result_out[28] ), .A2(_06081_ ), .B1(_06082_ ), .B2(_09378_ ), .ZN(_07916_ ) );
AOI21_X1 _22935_ ( .A(_06076_ ), .B1(_07915_ ), .B2(_07916_ ), .ZN(_00028_ ) );
OAI22_X1 _22936_ ( .A1(_09104_ ), .A2(_05731_ ), .B1(\u_gpr.gpr_wdata_$_ANDNOT__Y_30_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B2(_08928_ ), .ZN(_07917_ ) );
AND3_X1 _22937_ ( .A1(_06456_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06160_ ), .ZN(_07918_ ) );
AOI221_X4 _22938_ ( .A(_07918_ ), .B1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06923_ ), .C1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06176_ ), .ZN(_07919_ ) );
NAND3_X1 _22939_ ( .A1(_06152_ ), .A2(_06154_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07920_ ) );
NAND3_X1 _22940_ ( .A1(_07919_ ), .A2(_06368_ ), .A3(_07920_ ), .ZN(_07921_ ) );
AOI22_X1 _22941_ ( .A1(_06637_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06702_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07922_ ) );
OAI211_X1 _22942_ ( .A(_06798_ ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06600_ ), .C2(_06601_ ), .ZN(_07923_ ) );
NAND3_X1 _22943_ ( .A1(_06193_ ), .A2(_06194_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07924_ ) );
NAND3_X1 _22944_ ( .A1(_07922_ ), .A2(_07923_ ), .A3(_07924_ ), .ZN(_07925_ ) );
OAI211_X1 _22945_ ( .A(_07921_ ), .B(_06463_ ), .C1(_07008_ ), .C2(_07925_ ), .ZN(_07926_ ) );
AOI22_X1 _22946_ ( .A1(_06857_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06622_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07927_ ) );
OAI211_X1 _22947_ ( .A(_06798_ ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06353_ ), .C2(_06356_ ), .ZN(_07928_ ) );
NAND3_X1 _22948_ ( .A1(_06473_ ), .A2(_06515_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07929_ ) );
NAND4_X1 _22949_ ( .A1(_07927_ ), .A2(_06479_ ), .A3(_07928_ ), .A4(_07929_ ), .ZN(_07930_ ) );
AOI22_X1 _22950_ ( .A1(_06342_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06380_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07931_ ) );
OAI211_X1 _22951_ ( .A(_06931_ ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06353_ ), .C2(_06356_ ), .ZN(_07932_ ) );
NAND3_X1 _22952_ ( .A1(_06473_ ), .A2(_06515_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07933_ ) );
NAND4_X1 _22953_ ( .A1(_07931_ ), .A2(_06964_ ), .A3(_07932_ ), .A4(_07933_ ), .ZN(_07934_ ) );
NAND3_X1 _22954_ ( .A1(_10050_ ), .A2(_07930_ ), .A3(_07934_ ), .ZN(_07935_ ) );
AOI21_X1 _22955_ ( .A(_11196_ ), .B1(_07926_ ), .B2(_07935_ ), .ZN(_07936_ ) );
OAI211_X1 _22956_ ( .A(_06160_ ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06629_ ), .C2(_06630_ ), .ZN(_07937_ ) );
INV_X1 _22957_ ( .A(_07937_ ), .ZN(_07938_ ) );
AOI221_X4 _22958_ ( .A(_07938_ ), .B1(_06242_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .C2(_09627_ ), .ZN(_07939_ ) );
NAND3_X1 _22959_ ( .A1(_06625_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06783_ ), .ZN(_07940_ ) );
AOI21_X1 _22960_ ( .A(_06950_ ), .B1(_07939_ ), .B2(_07940_ ), .ZN(_07941_ ) );
AOI22_X1 _22961_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06522_ ), .B1(_07062_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07942_ ) );
AOI22_X1 _22962_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06638_ ), .B1(_06524_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07943_ ) );
AOI21_X1 _22963_ ( .A(_07031_ ), .B1(_07942_ ), .B2(_07943_ ), .ZN(_07944_ ) );
OAI21_X1 _22964_ ( .A(_06204_ ), .B1(_07941_ ), .B2(_07944_ ), .ZN(_07945_ ) );
AOI22_X1 _22965_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06205_ ), .B1(_06207_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07946_ ) );
AOI22_X1 _22966_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06211_ ), .B1(_06213_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07947_ ) );
NAND3_X1 _22967_ ( .A1(_07946_ ), .A2(_06209_ ), .A3(_07947_ ), .ZN(_07948_ ) );
AOI22_X1 _22968_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06216_ ), .B1(_06217_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07949_ ) );
AOI22_X1 _22969_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06220_ ), .B1(_06221_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07950_ ) );
NAND3_X1 _22970_ ( .A1(_07949_ ), .A2(_06219_ ), .A3(_07950_ ), .ZN(_07951_ ) );
NAND3_X1 _22971_ ( .A1(_06252_ ), .A2(_07948_ ), .A3(_07951_ ), .ZN(_07952_ ) );
AOI21_X1 _22972_ ( .A(_06186_ ), .B1(_07945_ ), .B2(_07952_ ), .ZN(_07953_ ) );
OAI21_X1 _22973_ ( .A(_10744_ ), .B1(_07936_ ), .B2(_07953_ ), .ZN(_07954_ ) );
AOI22_X1 _22974_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06365_ ), .B1(_06366_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07955_ ) );
AOI22_X1 _22975_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06369_ ), .B1(_06370_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07956_ ) );
NAND3_X1 _22976_ ( .A1(_07955_ ), .A2(_06368_ ), .A3(_07956_ ), .ZN(_07957_ ) );
AOI22_X1 _22977_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06637_ ), .B1(_06207_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07958_ ) );
AOI22_X1 _22978_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06794_ ), .B1(_06274_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07959_ ) );
NAND3_X1 _22979_ ( .A1(_07958_ ), .A2(_06329_ ), .A3(_07959_ ), .ZN(_07960_ ) );
NAND3_X1 _22980_ ( .A1(_06645_ ), .A2(_07957_ ), .A3(_07960_ ), .ZN(_07961_ ) );
AND3_X1 _22981_ ( .A1(_06440_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06598_ ), .ZN(_07962_ ) );
NAND3_X1 _22982_ ( .A1(_06434_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06436_ ), .ZN(_07963_ ) );
OAI211_X1 _22983_ ( .A(_06543_ ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06351_ ), .C2(_06354_ ), .ZN(_07964_ ) );
NAND2_X1 _22984_ ( .A1(_07963_ ), .A2(_07964_ ), .ZN(_07965_ ) );
AND3_X1 _22985_ ( .A1(_06434_ ), .A2(_06392_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07966_ ) );
NOR3_X1 _22986_ ( .A1(_07962_ ), .A2(_07965_ ), .A3(_07966_ ), .ZN(_07967_ ) );
AOI22_X1 _22987_ ( .A1(_06298_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06150_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07968_ ) );
NAND3_X1 _22988_ ( .A1(_07362_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06797_ ), .ZN(_07969_ ) );
NAND3_X1 _22989_ ( .A1(_06397_ ), .A2(_06598_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07970_ ) );
AND3_X1 _22990_ ( .A1(_07968_ ), .A2(_07969_ ), .A3(_07970_ ), .ZN(_07971_ ) );
MUX2_X1 _22991_ ( .A(_07967_ ), .B(_07971_ ), .S(_06158_ ), .Z(_07972_ ) );
OAI211_X1 _22992_ ( .A(_06654_ ), .B(_07961_ ), .C1(_07972_ ), .C2(_10261_ ), .ZN(_07973_ ) );
AOI22_X1 _22993_ ( .A1(_06593_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06322_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07974_ ) );
NAND3_X1 _22994_ ( .A1(_06459_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06311_ ), .ZN(_07975_ ) );
OAI211_X1 _22995_ ( .A(_06484_ ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06600_ ), .C2(_06601_ ), .ZN(_07976_ ) );
NAND4_X1 _22996_ ( .A1(_07974_ ), .A2(_06362_ ), .A3(_07975_ ), .A4(_07976_ ), .ZN(_07977_ ) );
AOI22_X1 _22997_ ( .A1(_06781_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06360_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07978_ ) );
NAND3_X1 _22998_ ( .A1(_06625_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06783_ ), .ZN(_07979_ ) );
OAI211_X1 _22999_ ( .A(_06484_ ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06600_ ), .C2(_06601_ ), .ZN(_07980_ ) );
NAND4_X1 _23000_ ( .A1(_07978_ ), .A2(_06565_ ), .A3(_07979_ ), .A4(_07980_ ), .ZN(_07981_ ) );
NAND3_X1 _23001_ ( .A1(_06573_ ), .A2(_07977_ ), .A3(_07981_ ), .ZN(_07982_ ) );
AOI22_X1 _23002_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06205_ ), .B1(_06217_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07983_ ) );
AOI22_X1 _23003_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06211_ ), .B1(_06274_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07984_ ) );
AOI21_X1 _23004_ ( .A(_06929_ ), .B1(_07983_ ), .B2(_07984_ ), .ZN(_07985_ ) );
AOI22_X1 _23005_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06382_ ), .B1(_06384_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_07986_ ) );
AOI22_X1 _23006_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06470_ ), .B1(_06425_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07987_ ) );
AOI21_X1 _23007_ ( .A(_06390_ ), .B1(_07986_ ), .B2(_07987_ ), .ZN(_07988_ ) );
OAI21_X1 _23008_ ( .A(_06252_ ), .B1(_07985_ ), .B2(_07988_ ), .ZN(_07989_ ) );
NAND3_X1 _23009_ ( .A1(_07982_ ), .A2(_09487_ ), .A3(_07989_ ), .ZN(_07990_ ) );
NAND3_X1 _23010_ ( .A1(_07973_ ), .A2(_06338_ ), .A3(_07990_ ), .ZN(_07991_ ) );
AOI21_X1 _23011_ ( .A(_02457_ ), .B1(_07954_ ), .B2(_07991_ ), .ZN(_07992_ ) );
AND3_X1 _23012_ ( .A1(_10430_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06391_ ), .ZN(_07993_ ) );
AOI221_X4 _23013_ ( .A(_07993_ ), .B1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06430_ ), .C1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C2(_06206_ ), .ZN(_07994_ ) );
NAND3_X1 _23014_ ( .A1(_09071_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06675_ ), .ZN(_07995_ ) );
NAND3_X1 _23015_ ( .A1(_07994_ ), .A2(_06300_ ), .A3(_07995_ ), .ZN(_07996_ ) );
AOI22_X1 _23016_ ( .A1(_06593_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06306_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07997_ ) );
NAND3_X1 _23017_ ( .A1(_06309_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06590_ ), .ZN(_07998_ ) );
NAND3_X1 _23018_ ( .A1(_06246_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06311_ ), .ZN(_07999_ ) );
NAND4_X1 _23019_ ( .A1(_07997_ ), .A2(_06308_ ), .A3(_07998_ ), .A4(_07999_ ), .ZN(_08000_ ) );
NAND3_X1 _23020_ ( .A1(_07996_ ), .A2(_06303_ ), .A3(_08000_ ), .ZN(_08001_ ) );
AOI22_X1 _23021_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06316_ ), .B1(_06318_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08002_ ) );
AOI22_X1 _23022_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06321_ ), .B1(_06322_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08003_ ) );
NAND3_X1 _23023_ ( .A1(_08002_ ), .A2(_06320_ ), .A3(_08003_ ), .ZN(_08004_ ) );
AOI22_X1 _23024_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06757_ ), .B1(_06306_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08005_ ) );
AOI22_X1 _23025_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06365_ ), .B1(_06263_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08006_ ) );
NAND3_X1 _23026_ ( .A1(_08005_ ), .A2(_06611_ ), .A3(_08006_ ), .ZN(_08007_ ) );
NAND3_X1 _23027_ ( .A1(_06315_ ), .A2(_08004_ ), .A3(_08007_ ), .ZN(_08008_ ) );
NAND3_X1 _23028_ ( .A1(_08001_ ), .A2(_11056_ ), .A3(_08008_ ), .ZN(_08009_ ) );
AOI22_X1 _23029_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06697_ ), .B1(_06360_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08010_ ) );
NAND3_X1 _23030_ ( .A1(_06625_ ), .A2(_06331_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08011_ ) );
NAND3_X1 _23031_ ( .A1(_06330_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06783_ ), .ZN(_08012_ ) );
NAND4_X1 _23032_ ( .A1(_08010_ ), .A2(_06565_ ), .A3(_08011_ ), .A4(_08012_ ), .ZN(_08013_ ) );
AOI22_X1 _23033_ ( .A1(_06346_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06327_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08014_ ) );
NAND3_X1 _23034_ ( .A1(_06330_ ), .A2(_06331_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08015_ ) );
OAI211_X1 _23035_ ( .A(_06798_ ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06353_ ), .C2(_06356_ ), .ZN(_08016_ ) );
NAND4_X1 _23036_ ( .A1(_08014_ ), .A2(_06219_ ), .A3(_08015_ ), .A4(_08016_ ), .ZN(_08017_ ) );
NAND3_X1 _23037_ ( .A1(_06315_ ), .A2(_08013_ ), .A3(_08017_ ), .ZN(_08018_ ) );
AOI22_X1 _23038_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06342_ ), .B1(_06343_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08019_ ) );
AOI22_X1 _23039_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06594_ ), .B1(_06380_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08020_ ) );
NAND3_X1 _23040_ ( .A1(_08019_ ), .A2(_06368_ ), .A3(_08020_ ), .ZN(_08021_ ) );
AOI22_X1 _23041_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06794_ ), .B1(_06702_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08022_ ) );
NAND3_X1 _23042_ ( .A1(_06483_ ), .A2(_06599_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08023_ ) );
NAND3_X1 _23043_ ( .A1(_06166_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06798_ ), .ZN(_08024_ ) );
NAND4_X1 _23044_ ( .A1(_08022_ ), .A2(_06514_ ), .A3(_08023_ ), .A4(_08024_ ), .ZN(_08025_ ) );
NAND3_X1 _23045_ ( .A1(_09056_ ), .A2(_08021_ ), .A3(_08025_ ), .ZN(_08026_ ) );
NAND3_X1 _23046_ ( .A1(_08018_ ), .A2(_09487_ ), .A3(_08026_ ), .ZN(_08027_ ) );
NAND3_X1 _23047_ ( .A1(_08009_ ), .A2(_06338_ ), .A3(_08027_ ), .ZN(_08028_ ) );
AOI22_X1 _23048_ ( .A1(_06836_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06221_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08029_ ) );
OAI211_X1 _23049_ ( .A(_06408_ ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06480_ ), .C2(_06481_ ), .ZN(_08030_ ) );
NAND3_X1 _23050_ ( .A1(_06492_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06931_ ), .ZN(_08031_ ) );
NAND4_X1 _23051_ ( .A1(_08029_ ), .A2(_06973_ ), .A3(_08030_ ), .A4(_08031_ ), .ZN(_08032_ ) );
AOI22_X1 _23052_ ( .A1(_06421_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06422_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_08033_ ) );
NAND3_X1 _23053_ ( .A1(_06492_ ), .A2(_06167_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08034_ ) );
OAI211_X1 _23054_ ( .A(_06978_ ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06394_ ), .C2(_06395_ ), .ZN(_08035_ ) );
NAND4_X1 _23055_ ( .A1(_08033_ ), .A2(_06255_ ), .A3(_08034_ ), .A4(_08035_ ), .ZN(_08036_ ) );
NAND3_X1 _23056_ ( .A1(_06254_ ), .A2(_08032_ ), .A3(_08036_ ), .ZN(_08037_ ) );
AOI22_X1 _23057_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06794_ ), .B1(_06274_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08038_ ) );
AOI22_X1 _23058_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06267_ ), .B1(_09795_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08039_ ) );
NAND3_X1 _23059_ ( .A1(_08038_ ), .A2(_06700_ ), .A3(_08039_ ), .ZN(_08040_ ) );
AOI22_X1 _23060_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06382_ ), .B1(_06540_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08041_ ) );
AOI22_X1 _23061_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06477_ ), .B1(_06425_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08042_ ) );
NAND3_X1 _23062_ ( .A1(_08041_ ), .A2(_06514_ ), .A3(_08042_ ), .ZN(_08043_ ) );
NAND3_X1 _23063_ ( .A1(_06388_ ), .A2(_08040_ ), .A3(_08043_ ), .ZN(_08044_ ) );
AOI21_X1 _23064_ ( .A(_06186_ ), .B1(_08037_ ), .B2(_08044_ ), .ZN(_08045_ ) );
AOI22_X1 _23065_ ( .A1(_06207_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06524_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08046_ ) );
NAND3_X1 _23066_ ( .A1(_06407_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06401_ ), .ZN(_08047_ ) );
OAI211_X1 _23067_ ( .A(_06544_ ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06417_ ), .C2(_06418_ ), .ZN(_08048_ ) );
NAND4_X1 _23068_ ( .A1(_08046_ ), .A2(_06390_ ), .A3(_08047_ ), .A4(_08048_ ), .ZN(_08049_ ) );
AOI22_X1 _23069_ ( .A1(_07061_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06288_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_08050_ ) );
NAND3_X1 _23070_ ( .A1(_06407_ ), .A2(_06939_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08051_ ) );
OAI211_X1 _23071_ ( .A(_09094_ ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06417_ ), .C2(_06418_ ), .ZN(_08052_ ) );
NAND4_X1 _23072_ ( .A1(_08050_ ), .A2(_07031_ ), .A3(_08051_ ), .A4(_08052_ ), .ZN(_08053_ ) );
NAND3_X1 _23073_ ( .A1(_06414_ ), .A2(_08049_ ), .A3(_08053_ ), .ZN(_08054_ ) );
AOI22_X1 _23074_ ( .A1(_06429_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06431_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_08055_ ) );
NAND3_X1 _23075_ ( .A1(_06435_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06437_ ), .ZN(_08056_ ) );
NAND3_X1 _23076_ ( .A1(_06441_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06393_ ), .ZN(_08057_ ) );
NAND4_X1 _23077_ ( .A1(_08055_ ), .A2(_06433_ ), .A3(_08056_ ), .A4(_08057_ ), .ZN(_08058_ ) );
AOI22_X1 _23078_ ( .A1(_06286_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06445_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08059_ ) );
NAND3_X1 _23079_ ( .A1(_06435_ ), .A2(_06393_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08060_ ) );
NAND3_X1 _23080_ ( .A1(_06448_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06544_ ), .ZN(_08061_ ) );
NAND4_X1 _23081_ ( .A1(_08059_ ), .A2(_06197_ ), .A3(_08060_ ), .A4(_08061_ ), .ZN(_08062_ ) );
NAND3_X1 _23082_ ( .A1(_06500_ ), .A2(_08058_ ), .A3(_08062_ ), .ZN(_08063_ ) );
AOI21_X1 _23083_ ( .A(_06413_ ), .B1(_08054_ ), .B2(_08063_ ), .ZN(_08064_ ) );
OAI21_X1 _23084_ ( .A(_06227_ ), .B1(_08045_ ), .B2(_08064_ ), .ZN(_08065_ ) );
AOI21_X1 _23085_ ( .A(_09604_ ), .B1(_08028_ ), .B2(_08065_ ), .ZN(_08066_ ) );
OAI21_X1 _23086_ ( .A(_09138_ ), .B1(_07992_ ), .B2(_08066_ ), .ZN(_08067_ ) );
NAND3_X1 _23087_ ( .A1(_06145_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06296_ ), .ZN(_08068_ ) );
INV_X1 _23088_ ( .A(_08068_ ), .ZN(_08069_ ) );
AOI221_X4 _23089_ ( .A(_08069_ ), .B1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06149_ ), .C1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06424_ ), .ZN(_08070_ ) );
NAND3_X1 _23090_ ( .A1(_06568_ ), .A2(_06569_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08071_ ) );
AOI21_X1 _23091_ ( .A(_06209_ ), .B1(_08070_ ), .B2(_08071_ ), .ZN(_08072_ ) );
OAI211_X1 _23092_ ( .A(_06187_ ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06629_ ), .C2(_06630_ ), .ZN(_08073_ ) );
INV_X1 _23093_ ( .A(_08073_ ), .ZN(_08074_ ) );
AOI221_X4 _23094_ ( .A(_08074_ ), .B1(_06923_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06190_ ), .ZN(_08075_ ) );
NAND3_X1 _23095_ ( .A1(_06193_ ), .A2(_06194_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08076_ ) );
AOI21_X1 _23096_ ( .A(_06405_ ), .B1(_08075_ ), .B2(_08076_ ), .ZN(_08077_ ) );
NOR3_X1 _23097_ ( .A1(_08072_ ), .A2(_08077_ ), .A3(_06388_ ), .ZN(_08078_ ) );
AOI22_X1 _23098_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06177_ ), .B1(_06181_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08079_ ) );
AOI22_X1 _23099_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06288_ ), .B1(_06289_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08080_ ) );
AOI21_X1 _23100_ ( .A(_06495_ ), .B1(_08079_ ), .B2(_08080_ ), .ZN(_08081_ ) );
AOI22_X1 _23101_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06304_ ), .B1(_06504_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08082_ ) );
AOI22_X1 _23102_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06179_ ), .B1(_06506_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08083_ ) );
AOI21_X1 _23103_ ( .A(_06244_ ), .B1(_08082_ ), .B2(_08083_ ), .ZN(_08084_ ) );
NOR3_X1 _23104_ ( .A1(_06414_ ), .A2(_08081_ ), .A3(_08084_ ), .ZN(_08085_ ) );
NOR3_X1 _23105_ ( .A1(_08078_ ), .A2(_06654_ ), .A3(_08085_ ), .ZN(_08086_ ) );
AND3_X1 _23106_ ( .A1(_06159_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06187_ ), .ZN(_08087_ ) );
AOI221_X4 _23107_ ( .A(_08087_ ), .B1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06189_ ), .C1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .C2(_09627_ ), .ZN(_08088_ ) );
NAND3_X1 _23108_ ( .A1(_06246_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06311_ ), .ZN(_08089_ ) );
NAND3_X1 _23109_ ( .A1(_08088_ ), .A2(_06329_ ), .A3(_08089_ ), .ZN(_08090_ ) );
MUX2_X1 _23110_ ( .A(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .S(_06199_ ), .Z(_08091_ ) );
MUX2_X1 _23111_ ( .A(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .S(_06464_ ), .Z(_08092_ ) );
MUX2_X1 _23112_ ( .A(_08091_ ), .B(_08092_ ), .S(_06448_ ), .Z(_08093_ ) );
OAI211_X1 _23113_ ( .A(_08090_ ), .B(_06388_ ), .C1(_06198_ ), .C2(_08093_ ), .ZN(_08094_ ) );
NAND3_X1 _23114_ ( .A1(_06671_ ), .A2(_09093_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08095_ ) );
INV_X1 _23115_ ( .A(_08095_ ), .ZN(_08096_ ) );
AOI221_X4 _23116_ ( .A(_08096_ ), .B1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06149_ ), .C1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06212_ ), .ZN(_08097_ ) );
NAND3_X1 _23117_ ( .A1(_06568_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06736_ ), .ZN(_08098_ ) );
NAND3_X1 _23118_ ( .A1(_08097_ ), .A2(_06611_ ), .A3(_08098_ ), .ZN(_08099_ ) );
OAI211_X1 _23119_ ( .A(_06256_ ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06629_ ), .C2(_06630_ ), .ZN(_08100_ ) );
INV_X1 _23120_ ( .A(_08100_ ), .ZN(_08101_ ) );
AOI221_X4 _23121_ ( .A(_08101_ ), .B1(_06231_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06176_ ), .ZN(_08102_ ) );
NAND3_X1 _23122_ ( .A1(_06152_ ), .A2(_06154_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08103_ ) );
NAND3_X1 _23123_ ( .A1(_08102_ ), .A2(_06368_ ), .A3(_08103_ ), .ZN(_08104_ ) );
NAND3_X1 _23124_ ( .A1(_08099_ ), .A2(_06204_ ), .A3(_08104_ ), .ZN(_08105_ ) );
AOI21_X1 _23125_ ( .A(_09594_ ), .B1(_08094_ ), .B2(_08105_ ), .ZN(_08106_ ) );
OAI21_X1 _23126_ ( .A(_06143_ ), .B1(_08086_ ), .B2(_08106_ ), .ZN(_08107_ ) );
NAND3_X1 _23127_ ( .A1(_06671_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06399_ ), .ZN(_08108_ ) );
INV_X1 _23128_ ( .A(_08108_ ), .ZN(_08109_ ) );
AOI221_X4 _23129_ ( .A(_08109_ ), .B1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06430_ ), .C1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06326_ ), .ZN(_08110_ ) );
NAND3_X1 _23130_ ( .A1(_06561_ ), .A2(_06562_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08111_ ) );
NAND3_X1 _23131_ ( .A1(_08110_ ), .A2(_06576_ ), .A3(_08111_ ), .ZN(_08112_ ) );
OAI211_X1 _23132_ ( .A(_06678_ ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06629_ ), .C2(_06630_ ), .ZN(_08113_ ) );
INV_X1 _23133_ ( .A(_08113_ ), .ZN(_08114_ ) );
AOI221_X4 _23134_ ( .A(_08114_ ), .B1(_06716_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06285_ ), .ZN(_08115_ ) );
NAND3_X1 _23135_ ( .A1(_06568_ ), .A2(_06569_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08116_ ) );
NAND3_X1 _23136_ ( .A1(_08115_ ), .A2(_06245_ ), .A3(_08116_ ), .ZN(_08117_ ) );
NAND3_X1 _23137_ ( .A1(_08112_ ), .A2(_06890_ ), .A3(_08117_ ), .ZN(_08118_ ) );
AOI22_X1 _23138_ ( .A1(_06317_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06212_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08119_ ) );
NAND3_X1 _23139_ ( .A1(_06165_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06797_ ), .ZN(_08120_ ) );
NAND3_X1 _23140_ ( .A1(_07362_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06797_ ), .ZN(_08121_ ) );
AND3_X1 _23141_ ( .A1(_08119_ ), .A2(_08120_ ), .A3(_08121_ ), .ZN(_08122_ ) );
AOI22_X1 _23142_ ( .A1(_06317_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06212_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08123_ ) );
NAND3_X1 _23143_ ( .A1(_06165_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06248_ ), .ZN(_08124_ ) );
NAND3_X1 _23144_ ( .A1(_07362_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06797_ ), .ZN(_08125_ ) );
AND3_X1 _23145_ ( .A1(_08123_ ), .A2(_08124_ ), .A3(_08125_ ), .ZN(_08126_ ) );
MUX2_X1 _23146_ ( .A(_08122_ ), .B(_08126_ ), .S(_06405_ ), .Z(_08127_ ) );
OAI211_X1 _23147_ ( .A(_08118_ ), .B(_09487_ ), .C1(_08127_ ), .C2(_10261_ ), .ZN(_08128_ ) );
AOI22_X1 _23148_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06574_ ), .B1(_06781_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08129_ ) );
AOI22_X1 _23149_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06339_ ), .B1(_09530_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08130_ ) );
NAND3_X1 _23150_ ( .A1(_08129_ ), .A2(_06300_ ), .A3(_08130_ ), .ZN(_08131_ ) );
AOI22_X1 _23151_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06574_ ), .B1(_06781_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08132_ ) );
AOI22_X1 _23152_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06339_ ), .B1(_06340_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08133_ ) );
NAND3_X1 _23153_ ( .A1(_08132_ ), .A2(_06576_ ), .A3(_08133_ ), .ZN(_08134_ ) );
NAND3_X1 _23154_ ( .A1(_10261_ ), .A2(_08131_ ), .A3(_08134_ ), .ZN(_08135_ ) );
AOI22_X1 _23155_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06316_ ), .B1(_06476_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08136_ ) );
AOI22_X1 _23156_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06757_ ), .B1(_06322_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08137_ ) );
NAND3_X1 _23157_ ( .A1(_08136_ ), .A2(_06582_ ), .A3(_08137_ ), .ZN(_08138_ ) );
AOI22_X1 _23158_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06316_ ), .B1(_06318_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08139_ ) );
AOI22_X1 _23159_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06321_ ), .B1(_06322_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08140_ ) );
NAND3_X1 _23160_ ( .A1(_08139_ ), .A2(_06234_ ), .A3(_08140_ ), .ZN(_08141_ ) );
NAND3_X1 _23161_ ( .A1(_06303_ ), .A2(_08138_ ), .A3(_08141_ ), .ZN(_08142_ ) );
NAND3_X1 _23162_ ( .A1(_08135_ ), .A2(_11056_ ), .A3(_08142_ ), .ZN(_08143_ ) );
NAND3_X1 _23163_ ( .A1(_08128_ ), .A2(_10744_ ), .A3(_08143_ ), .ZN(_08144_ ) );
NAND3_X1 _23164_ ( .A1(_08107_ ), .A2(_08144_ ), .A3(_09604_ ), .ZN(_08145_ ) );
AND3_X1 _23165_ ( .A1(_06439_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06146_ ), .ZN(_08146_ ) );
AOI221_X4 _23166_ ( .A(_08146_ ), .B1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06716_ ), .C1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06298_ ), .ZN(_08147_ ) );
NAND3_X1 _23167_ ( .A1(_06718_ ), .A2(_09095_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08148_ ) );
NAND3_X1 _23168_ ( .A1(_08147_ ), .A2(_06576_ ), .A3(_08148_ ), .ZN(_08149_ ) );
AND3_X1 _23169_ ( .A1(_06557_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06678_ ), .ZN(_08150_ ) );
AOI221_X4 _23170_ ( .A(_08150_ ), .B1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06559_ ), .C1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06232_ ), .ZN(_08151_ ) );
NAND3_X1 _23171_ ( .A1(_06235_ ), .A2(_06236_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08152_ ) );
NAND3_X1 _23172_ ( .A1(_08151_ ), .A2(_06582_ ), .A3(_08152_ ), .ZN(_08153_ ) );
NAND3_X1 _23173_ ( .A1(_08149_ ), .A2(_08153_ ), .A3(_10050_ ), .ZN(_08154_ ) );
AOI22_X1 _23174_ ( .A1(_06469_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06347_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_08155_ ) );
NAND3_X1 _23175_ ( .A1(_06330_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06783_ ), .ZN(_08156_ ) );
OAI211_X1 _23176_ ( .A(_06350_ ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(_06353_ ), .C2(_06356_ ), .ZN(_08157_ ) );
NAND4_X1 _23177_ ( .A1(_08155_ ), .A2(_06219_ ), .A3(_08156_ ), .A4(_08157_ ), .ZN(_08158_ ) );
AOI22_X1 _23178_ ( .A1(_06316_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_06369_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_08159_ ) );
AOI22_X1 _23179_ ( .A1(_06781_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_06327_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08160_ ) );
NAND3_X1 _23180_ ( .A1(_08159_ ), .A2(_08160_ ), .A3(_06596_ ), .ZN(_08161_ ) );
NAND3_X1 _23181_ ( .A1(_06890_ ), .A2(_08158_ ), .A3(_08161_ ), .ZN(_08162_ ) );
AOI21_X1 _23182_ ( .A(_11196_ ), .B1(_08154_ ), .B2(_08162_ ), .ZN(_08163_ ) );
NAND3_X1 _23183_ ( .A1(_06671_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06399_ ), .ZN(_08164_ ) );
INV_X1 _23184_ ( .A(_08164_ ), .ZN(_08165_ ) );
AOI221_X4 _23185_ ( .A(_08165_ ), .B1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06149_ ), .C1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06212_ ), .ZN(_08166_ ) );
NAND3_X1 _23186_ ( .A1(_06235_ ), .A2(_06236_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08167_ ) );
NAND3_X1 _23187_ ( .A1(_08166_ ), .A2(_06234_ ), .A3(_08167_ ), .ZN(_08168_ ) );
NAND3_X1 _23188_ ( .A1(_06145_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06296_ ), .ZN(_08169_ ) );
INV_X1 _23189_ ( .A(_08169_ ), .ZN(_08170_ ) );
AOI221_X4 _23190_ ( .A(_08170_ ), .B1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06149_ ), .C1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06424_ ), .ZN(_08171_ ) );
NAND3_X1 _23191_ ( .A1(_06925_ ), .A2(_06811_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08172_ ) );
NAND3_X1 _23192_ ( .A1(_08171_ ), .A2(_06596_ ), .A3(_08172_ ), .ZN(_08173_ ) );
NAND3_X1 _23193_ ( .A1(_08168_ ), .A2(_08173_ ), .A3(_06254_ ), .ZN(_08174_ ) );
AOI22_X1 _23194_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_09746_ ), .B1(_06540_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08175_ ) );
AOI22_X1 _23195_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06470_ ), .B1(_06864_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08176_ ) );
AOI21_X1 _23196_ ( .A(_06405_ ), .B1(_08175_ ), .B2(_08176_ ), .ZN(_08177_ ) );
AOI22_X1 _23197_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06444_ ), .B1(_06527_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08178_ ) );
AOI22_X1 _23198_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_09484_ ), .B1(_06268_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08179_ ) );
AOI21_X1 _23199_ ( .A(_06433_ ), .B1(_08178_ ), .B2(_08179_ ), .ZN(_08180_ ) );
OAI21_X1 _23200_ ( .A(_06684_ ), .B1(_08177_ ), .B2(_08180_ ), .ZN(_08181_ ) );
AOI21_X1 _23201_ ( .A(_06186_ ), .B1(_08174_ ), .B2(_08181_ ), .ZN(_08182_ ) );
OAI21_X1 _23202_ ( .A(_10744_ ), .B1(_08163_ ), .B2(_08182_ ), .ZN(_08183_ ) );
AND3_X1 _23203_ ( .A1(_06228_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A3(_06256_ ), .ZN(_08184_ ) );
AOI221_X4 _23204_ ( .A(_08184_ ), .B1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06242_ ), .C1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06285_ ), .ZN(_08185_ ) );
NAND3_X1 _23205_ ( .A1(_06619_ ), .A2(_06569_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08186_ ) );
NAND3_X1 _23206_ ( .A1(_08185_ ), .A2(_06245_ ), .A3(_08186_ ), .ZN(_08187_ ) );
MUX2_X1 _23207_ ( .A(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .S(_06464_ ), .Z(_08188_ ) );
MUX2_X1 _23208_ ( .A(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .S(_06722_ ), .Z(_08189_ ) );
MUX2_X1 _23209_ ( .A(_08188_ ), .B(_08189_ ), .S(_06448_ ), .Z(_08190_ ) );
OAI211_X1 _23210_ ( .A(_08187_ ), .B(_06645_ ), .C1(_07008_ ), .C2(_08190_ ), .ZN(_08191_ ) );
NAND3_X1 _23211_ ( .A1(_06145_ ), .A2(_06391_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08192_ ) );
INV_X1 _23212_ ( .A(_08192_ ), .ZN(_08193_ ) );
AOI221_X4 _23213_ ( .A(_08193_ ), .B1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06149_ ), .C1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C2(_06424_ ), .ZN(_08194_ ) );
NAND3_X1 _23214_ ( .A1(_06619_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06249_ ), .ZN(_08195_ ) );
AOI21_X1 _23215_ ( .A(_06479_ ), .B1(_08194_ ), .B2(_08195_ ), .ZN(_08196_ ) );
OAI211_X1 _23216_ ( .A(_06160_ ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06629_ ), .C2(_06630_ ), .ZN(_08197_ ) );
INV_X1 _23217_ ( .A(_08197_ ), .ZN(_08198_ ) );
AOI221_X4 _23218_ ( .A(_08198_ ), .B1(_06242_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .C2(_09627_ ), .ZN(_08199_ ) );
NAND3_X1 _23219_ ( .A1(_06625_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06783_ ), .ZN(_08200_ ) );
AOI21_X1 _23220_ ( .A(_06929_ ), .B1(_08199_ ), .B2(_08200_ ), .ZN(_08201_ ) );
OAI21_X1 _23221_ ( .A(_10050_ ), .B1(_08196_ ), .B2(_08201_ ), .ZN(_08202_ ) );
NAND3_X1 _23222_ ( .A1(_08191_ ), .A2(_10053_ ), .A3(_08202_ ), .ZN(_08203_ ) );
OAI211_X1 _23223_ ( .A(_06229_ ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06629_ ), .C2(_06630_ ), .ZN(_08204_ ) );
INV_X1 _23224_ ( .A(_08204_ ), .ZN(_08205_ ) );
AOI221_X4 _23225_ ( .A(_08205_ ), .B1(_06559_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .C2(_06176_ ), .ZN(_08206_ ) );
NAND3_X1 _23226_ ( .A1(_06925_ ), .A2(_06811_ ), .A3(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08207_ ) );
AOI21_X1 _23227_ ( .A(_06964_ ), .B1(_08206_ ), .B2(_08207_ ), .ZN(_08208_ ) );
OAI211_X1 _23228_ ( .A(_06160_ ), .B(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C1(_06629_ ), .C2(_06630_ ), .ZN(_08209_ ) );
INV_X1 _23229_ ( .A(_08209_ ), .ZN(_08210_ ) );
AOI221_X4 _23230_ ( .A(_08210_ ), .B1(_06923_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .C1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .C2(_09627_ ), .ZN(_08211_ ) );
NAND3_X1 _23231_ ( .A1(_06330_ ), .A2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A3(_06783_ ), .ZN(_08212_ ) );
AOI21_X1 _23232_ ( .A(_06950_ ), .B1(_08211_ ), .B2(_08212_ ), .ZN(_08213_ ) );
OAI21_X1 _23233_ ( .A(_06890_ ), .B1(_08208_ ), .B2(_08213_ ), .ZN(_08214_ ) );
AOI22_X1 _23234_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06205_ ), .B1(_06217_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08215_ ) );
AOI22_X1 _23235_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06211_ ), .B1(_06274_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08216_ ) );
AOI21_X1 _23236_ ( .A(_06929_ ), .B1(_08215_ ), .B2(_08216_ ), .ZN(_08217_ ) );
AOI22_X1 _23237_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .A2(_06382_ ), .B1(_06384_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_08218_ ) );
AOI22_X1 _23238_ ( .A1(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_06477_ ), .B1(_06425_ ), .B2(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08219_ ) );
AOI21_X1 _23239_ ( .A(_06390_ ), .B1(_08218_ ), .B2(_08219_ ), .ZN(_08220_ ) );
OAI21_X1 _23240_ ( .A(_06252_ ), .B1(_08217_ ), .B2(_08220_ ), .ZN(_08221_ ) );
NAND3_X1 _23241_ ( .A1(_08214_ ), .A2(_06654_ ), .A3(_08221_ ), .ZN(_08222_ ) );
NAND3_X1 _23242_ ( .A1(_08203_ ), .A2(_06338_ ), .A3(_08222_ ), .ZN(_08223_ ) );
NAND3_X1 _23243_ ( .A1(_08183_ ), .A2(_02457_ ), .A3(_08223_ ), .ZN(_08224_ ) );
NAND3_X1 _23244_ ( .A1(_08145_ ), .A2(_08224_ ), .A3(_09035_ ), .ZN(_08225_ ) );
AND3_X1 _23245_ ( .A1(_08067_ ), .A2(_08225_ ), .A3(_05734_ ), .ZN(\load_data_out[1] ) );
INV_X1 _23246_ ( .A(\load_data_out[1] ), .ZN(_08226_ ) );
OAI21_X1 _23247_ ( .A(_08226_ ), .B1(_09104_ ), .B2(_06130_ ), .ZN(_08227_ ) );
AOI21_X1 _23248_ ( .A(_07917_ ), .B1(_08227_ ), .B2(_06101_ ), .ZN(_08228_ ) );
NOR2_X1 _23249_ ( .A1(_08228_ ), .A2(_06137_ ), .ZN(_00029_ ) );
AND3_X1 _23250_ ( .A1(_10430_ ), .A2(\u_lsu.pmem[1696] ), .A3(_06722_ ), .ZN(_08229_ ) );
AOI221_X4 _23251_ ( .A(_08229_ ), .B1(\u_lsu.pmem[1664] ), .B2(_06506_ ), .C1(\u_lsu.pmem[1760] ), .C2(_09746_ ), .ZN(_08230_ ) );
BUF_X4 _23252_ ( .A(_09085_ ), .Z(_08231_ ) );
BUF_X4 _23253_ ( .A(_06718_ ), .Z(_08232_ ) );
BUF_X4 _23254_ ( .A(_06569_ ), .Z(_08233_ ) );
NAND3_X1 _23255_ ( .A1(_08232_ ), .A2(_08233_ ), .A3(\u_lsu.pmem[1728] ), .ZN(_08234_ ) );
NAND3_X1 _23256_ ( .A1(_08230_ ), .A2(_08231_ ), .A3(_08234_ ), .ZN(_08235_ ) );
BUF_X4 _23257_ ( .A(_06555_ ), .Z(_08236_ ) );
MUX2_X1 _23258_ ( .A(\u_lsu.pmem[1600] ), .B(\u_lsu.pmem[1632] ), .S(_06544_ ), .Z(_08237_ ) );
MUX2_X1 _23259_ ( .A(\u_lsu.pmem[1536] ), .B(\u_lsu.pmem[1568] ), .S(_06544_ ), .Z(_08238_ ) );
MUX2_X1 _23260_ ( .A(_08237_ ), .B(_08238_ ), .S(_10432_ ), .Z(_08239_ ) );
OAI211_X1 _23261_ ( .A(_08235_ ), .B(_08236_ ), .C1(\alu_result_out[4] ), .C2(_08239_ ), .ZN(_08240_ ) );
BUF_X2 _23262_ ( .A(_06245_ ), .Z(_08241_ ) );
BUF_X4 _23263_ ( .A(_06741_ ), .Z(_08242_ ) );
BUF_X4 _23264_ ( .A(_09530_ ), .Z(_08243_ ) );
AOI22_X1 _23265_ ( .A1(_08242_ ), .A2(\u_lsu.pmem[1856] ), .B1(_08243_ ), .B2(\u_lsu.pmem[1792] ), .ZN(_08244_ ) );
BUF_X4 _23266_ ( .A(_06736_ ), .Z(_08245_ ) );
OAI211_X1 _23267_ ( .A(_08245_ ), .B(\u_lsu.pmem[1824] ), .C1(_06743_ ), .C2(_06744_ ), .ZN(_08246_ ) );
BUF_X4 _23268_ ( .A(_09071_ ), .Z(_08247_ ) );
BUF_X2 _23269_ ( .A(_06736_ ), .Z(\alu_result_out[2] ) );
NAND3_X1 _23270_ ( .A1(_08247_ ), .A2(\u_lsu.pmem[1888] ), .A3(\alu_result_out[2] ), .ZN(_08248_ ) );
AND4_X1 _23271_ ( .A1(_08241_ ), .A2(_08244_ ), .A3(_08246_ ), .A4(_08248_ ), .ZN(_08249_ ) );
BUF_X4 _23272_ ( .A(_06304_ ), .Z(_08250_ ) );
BUF_X4 _23273_ ( .A(_08250_ ), .Z(_08251_ ) );
AOI22_X1 _23274_ ( .A1(_08251_ ), .A2(\u_lsu.pmem[2016] ), .B1(_08243_ ), .B2(\u_lsu.pmem[1920] ), .ZN(_08252_ ) );
OAI211_X1 _23275_ ( .A(_08245_ ), .B(\u_lsu.pmem[1952] ), .C1(_06743_ ), .C2(_06744_ ), .ZN(_08253_ ) );
NAND3_X1 _23276_ ( .A1(_08232_ ), .A2(_08233_ ), .A3(\u_lsu.pmem[1984] ), .ZN(_08254_ ) );
NAND4_X1 _23277_ ( .A1(_08252_ ), .A2(_08231_ ), .A3(_08253_ ), .A4(_08254_ ), .ZN(_08255_ ) );
NAND2_X1 _23278_ ( .A1(_10529_ ), .A2(_08255_ ), .ZN(_08256_ ) );
OAI211_X1 _23279_ ( .A(_08240_ ), .B(_09784_ ), .C1(_08249_ ), .C2(_08256_ ), .ZN(_08257_ ) );
AOI22_X1 _23280_ ( .A1(\u_lsu.pmem[1056] ), .A2(_06697_ ), .B1(_06327_ ), .B2(\u_lsu.pmem[1024] ), .ZN(_08258_ ) );
NAND3_X1 _23281_ ( .A1(_06309_ ), .A2(\u_lsu.pmem[1120] ), .A3(_06590_ ), .ZN(_08259_ ) );
NAND3_X1 _23282_ ( .A1(_06459_ ), .A2(_06460_ ), .A3(\u_lsu.pmem[1088] ), .ZN(_08260_ ) );
NAND3_X1 _23283_ ( .A1(_08258_ ), .A2(_08259_ ), .A3(_08260_ ), .ZN(_08261_ ) );
AOI22_X1 _23284_ ( .A1(\u_lsu.pmem[1184] ), .A2(_06697_ ), .B1(_06360_ ), .B2(\u_lsu.pmem[1152] ), .ZN(_08262_ ) );
NAND3_X1 _23285_ ( .A1(_06925_ ), .A2(_06811_ ), .A3(\u_lsu.pmem[1216] ), .ZN(_08263_ ) );
NAND3_X1 _23286_ ( .A1(_06152_ ), .A2(\u_lsu.pmem[1248] ), .A3(_06590_ ), .ZN(_08264_ ) );
NAND3_X1 _23287_ ( .A1(_08262_ ), .A2(_08263_ ), .A3(_08264_ ), .ZN(_08265_ ) );
MUX2_X1 _23288_ ( .A(_08261_ ), .B(_08265_ ), .S(_09085_ ), .Z(_08266_ ) );
AOI22_X1 _23289_ ( .A1(\u_lsu.pmem[1312] ), .A2(_06697_ ), .B1(_06360_ ), .B2(\u_lsu.pmem[1280] ), .ZN(_08267_ ) );
NAND3_X1 _23290_ ( .A1(_06925_ ), .A2(\u_lsu.pmem[1376] ), .A3(_06249_ ), .ZN(_08268_ ) );
NAND3_X1 _23291_ ( .A1(_06152_ ), .A2(_06154_ ), .A3(\u_lsu.pmem[1344] ), .ZN(_08269_ ) );
NAND3_X1 _23292_ ( .A1(_08267_ ), .A2(_08268_ ), .A3(_08269_ ), .ZN(_08270_ ) );
AOI22_X1 _23293_ ( .A1(\u_lsu.pmem[1504] ), .A2(_06605_ ), .B1(_06318_ ), .B2(\u_lsu.pmem[1472] ), .ZN(_08271_ ) );
AOI22_X1 _23294_ ( .A1(\u_lsu.pmem[1440] ), .A2(_06757_ ), .B1(_06322_ ), .B2(\u_lsu.pmem[1408] ), .ZN(_08272_ ) );
NAND2_X1 _23295_ ( .A1(_08271_ ), .A2(_08272_ ), .ZN(_08273_ ) );
MUX2_X1 _23296_ ( .A(_08270_ ), .B(_08273_ ), .S(_09085_ ), .Z(_08274_ ) );
MUX2_X1 _23297_ ( .A(_08266_ ), .B(_08274_ ), .S(_10529_ ), .Z(_08275_ ) );
OAI211_X1 _23298_ ( .A(_08257_ ), .B(_10286_ ), .C1(_08275_ ), .C2(_09785_ ), .ZN(_08276_ ) );
AND3_X1 _23299_ ( .A1(_10430_ ), .A2(\u_lsu.pmem[32] ), .A3(_06436_ ), .ZN(_08277_ ) );
AOI221_X4 _23300_ ( .A(_08277_ ), .B1(\u_lsu.pmem[0] ), .B2(_06915_ ), .C1(\u_lsu.pmem[64] ), .C2(_06781_ ), .ZN(_08278_ ) );
NAND3_X1 _23301_ ( .A1(\alu_result_out[3] ), .A2(\u_lsu.pmem[96] ), .A3(\alu_result_out[2] ), .ZN(_08279_ ) );
AOI21_X1 _23302_ ( .A(_08231_ ), .B1(_08278_ ), .B2(_08279_ ), .ZN(_08280_ ) );
AND3_X1 _23303_ ( .A1(_10430_ ), .A2(\u_lsu.pmem[160] ), .A3(_06543_ ), .ZN(_08281_ ) );
AOI221_X4 _23304_ ( .A(_08281_ ), .B1(\u_lsu.pmem[128] ), .B2(_06289_ ), .C1(\u_lsu.pmem[224] ), .C2(_06205_ ), .ZN(_08282_ ) );
BUF_X4 _23305_ ( .A(_09095_ ), .Z(_08283_ ) );
NAND3_X1 _23306_ ( .A1(_08247_ ), .A2(_08283_ ), .A3(\u_lsu.pmem[192] ), .ZN(_08284_ ) );
AOI21_X1 _23307_ ( .A(_07008_ ), .B1(_08282_ ), .B2(_08284_ ), .ZN(_08285_ ) );
OAI21_X1 _23308_ ( .A(_09888_ ), .B1(_08280_ ), .B2(_08285_ ), .ZN(_08286_ ) );
AND3_X1 _23309_ ( .A1(_10432_ ), .A2(\u_lsu.pmem[256] ), .A3(_06569_ ), .ZN(_08287_ ) );
NAND3_X1 _23310_ ( .A1(_06459_ ), .A2(\u_lsu.pmem[352] ), .A3(_06311_ ), .ZN(_08288_ ) );
OAI211_X1 _23311_ ( .A(_06484_ ), .B(\u_lsu.pmem[288] ), .C1(_06600_ ), .C2(_06601_ ), .ZN(_08289_ ) );
NAND2_X1 _23312_ ( .A1(_08288_ ), .A2(_08289_ ), .ZN(_08290_ ) );
AND3_X1 _23313_ ( .A1(_06483_ ), .A2(_06599_ ), .A3(\u_lsu.pmem[320] ), .ZN(_08291_ ) );
NOR3_X1 _23314_ ( .A1(_08287_ ), .A2(_08290_ ), .A3(_08291_ ), .ZN(_08292_ ) );
AND3_X1 _23315_ ( .A1(_10432_ ), .A2(\u_lsu.pmem[384] ), .A3(_06569_ ), .ZN(_08293_ ) );
NAND3_X1 _23316_ ( .A1(_06459_ ), .A2(_06460_ ), .A3(\u_lsu.pmem[448] ), .ZN(_08294_ ) );
OAI211_X1 _23317_ ( .A(_06484_ ), .B(\u_lsu.pmem[416] ), .C1(_06600_ ), .C2(_06601_ ), .ZN(_08295_ ) );
NAND2_X1 _23318_ ( .A1(_08294_ ), .A2(_08295_ ), .ZN(_08296_ ) );
AND3_X1 _23319_ ( .A1(_06483_ ), .A2(\u_lsu.pmem[480] ), .A3(_06484_ ), .ZN(_08297_ ) );
NOR3_X1 _23320_ ( .A1(_08293_ ), .A2(_08296_ ), .A3(_08297_ ), .ZN(_08298_ ) );
MUX2_X1 _23321_ ( .A(_08292_ ), .B(_08298_ ), .S(_06721_ ), .Z(_08299_ ) );
OAI211_X1 _23322_ ( .A(_08286_ ), .B(_09666_ ), .C1(_09888_ ), .C2(_08299_ ), .ZN(_08300_ ) );
AND3_X1 _23323_ ( .A1(_07362_ ), .A2(\u_lsu.pmem[800] ), .A3(_06797_ ), .ZN(_08301_ ) );
AOI221_X4 _23324_ ( .A(_08301_ ), .B1(\u_lsu.pmem[768] ), .B2(_06322_ ), .C1(\u_lsu.pmem[864] ), .C2(_08250_ ), .ZN(_08302_ ) );
NAND3_X1 _23325_ ( .A1(\alu_result_out[3] ), .A2(_09096_ ), .A3(\u_lsu.pmem[832] ), .ZN(_08303_ ) );
NAND3_X1 _23326_ ( .A1(_08302_ ), .A2(_07009_ ), .A3(_08303_ ), .ZN(_08304_ ) );
AND3_X1 _23327_ ( .A1(_07362_ ), .A2(\u_lsu.pmem[928] ), .A3(_06797_ ), .ZN(_08305_ ) );
AOI221_X4 _23328_ ( .A(_08305_ ), .B1(\u_lsu.pmem[896] ), .B2(_06622_ ), .C1(\u_lsu.pmem[992] ), .C2(_08250_ ), .ZN(_08306_ ) );
NAND3_X1 _23329_ ( .A1(\alu_result_out[3] ), .A2(_09096_ ), .A3(\u_lsu.pmem[960] ), .ZN(_08307_ ) );
NAND3_X1 _23330_ ( .A1(_08306_ ), .A2(\alu_result_out[4] ), .A3(_08307_ ), .ZN(_08308_ ) );
NAND3_X1 _23331_ ( .A1(_08304_ ), .A2(_08308_ ), .A3(\alu_result_out[5] ), .ZN(_08309_ ) );
AND3_X1 _23332_ ( .A1(_06434_ ), .A2(_06392_ ), .A3(\u_lsu.pmem[704] ), .ZN(_08310_ ) );
AOI221_X4 _23333_ ( .A(_08310_ ), .B1(\u_lsu.pmem[640] ), .B2(_06915_ ), .C1(\u_lsu.pmem[736] ), .C2(_06346_ ), .ZN(_08311_ ) );
BUF_X4 _23334_ ( .A(_09085_ ), .Z(_08312_ ) );
NAND3_X1 _23335_ ( .A1(_10433_ ), .A2(\u_lsu.pmem[672] ), .A3(\alu_result_out[2] ), .ZN(_08313_ ) );
NAND3_X1 _23336_ ( .A1(_08311_ ), .A2(_08312_ ), .A3(_08313_ ), .ZN(_08314_ ) );
MUX2_X1 _23337_ ( .A(\u_lsu.pmem[576] ), .B(\u_lsu.pmem[608] ), .S(_06437_ ), .Z(_08315_ ) );
MUX2_X1 _23338_ ( .A(\u_lsu.pmem[512] ), .B(\u_lsu.pmem[544] ), .S(_06437_ ), .Z(_08316_ ) );
MUX2_X1 _23339_ ( .A(_08315_ ), .B(_08316_ ), .S(_10432_ ), .Z(_08317_ ) );
OAI211_X1 _23340_ ( .A(_08314_ ), .B(_08236_ ), .C1(\alu_result_out[4] ), .C2(_08317_ ), .ZN(_08318_ ) );
NAND3_X1 _23341_ ( .A1(_08309_ ), .A2(_09785_ ), .A3(_08318_ ), .ZN(_08319_ ) );
NAND3_X1 _23342_ ( .A1(_08300_ ), .A2(_08319_ ), .A3(_09805_ ), .ZN(_08320_ ) );
NAND3_X1 _23343_ ( .A1(_08276_ ), .A2(_08320_ ), .A3(_02484_ ), .ZN(_08321_ ) );
AND3_X1 _23344_ ( .A1(_06440_ ), .A2(\u_lsu.pmem[2848] ), .A3(_06400_ ), .ZN(_08322_ ) );
AOI221_X4 _23345_ ( .A(_08322_ ), .B1(\u_lsu.pmem[2816] ), .B2(_06213_ ), .C1(\u_lsu.pmem[2912] ), .C2(_06305_ ), .ZN(_08323_ ) );
NAND3_X1 _23346_ ( .A1(\alu_result_out[3] ), .A2(_09096_ ), .A3(\u_lsu.pmem[2880] ), .ZN(_08324_ ) );
NAND3_X1 _23347_ ( .A1(_08323_ ), .A2(_07009_ ), .A3(_08324_ ), .ZN(_08325_ ) );
MUX2_X1 _23348_ ( .A(\u_lsu.pmem[3008] ), .B(\u_lsu.pmem[3040] ), .S(_06401_ ), .Z(_08326_ ) );
MUX2_X1 _23349_ ( .A(\u_lsu.pmem[2944] ), .B(\u_lsu.pmem[2976] ), .S(_06401_ ), .Z(_08327_ ) );
MUX2_X1 _23350_ ( .A(_08326_ ), .B(_08327_ ), .S(_10433_ ), .Z(_08328_ ) );
OAI211_X1 _23351_ ( .A(_08325_ ), .B(_10529_ ), .C1(_07009_ ), .C2(_08328_ ), .ZN(_08329_ ) );
BUF_X4 _23352_ ( .A(_08250_ ), .Z(_08330_ ) );
BUF_X4 _23353_ ( .A(_06339_ ), .Z(_08331_ ) );
AOI22_X1 _23354_ ( .A1(_08330_ ), .A2(\u_lsu.pmem[2656] ), .B1(_08331_ ), .B2(\u_lsu.pmem[2592] ), .ZN(_08332_ ) );
OAI211_X1 _23355_ ( .A(_08283_ ), .B(\u_lsu.pmem[2560] ), .C1(_06743_ ), .C2(_06744_ ), .ZN(_08333_ ) );
NAND3_X1 _23356_ ( .A1(_08247_ ), .A2(_08283_ ), .A3(\u_lsu.pmem[2624] ), .ZN(_08334_ ) );
NAND4_X1 _23357_ ( .A1(_08332_ ), .A2(_07009_ ), .A3(_08333_ ), .A4(_08334_ ), .ZN(_08335_ ) );
BUF_X4 _23358_ ( .A(_06339_ ), .Z(_08336_ ) );
AOI22_X1 _23359_ ( .A1(_08242_ ), .A2(\u_lsu.pmem[2752] ), .B1(_08336_ ), .B2(\u_lsu.pmem[2720] ), .ZN(_08337_ ) );
OAI211_X1 _23360_ ( .A(_08283_ ), .B(\u_lsu.pmem[2688] ), .C1(_06743_ ), .C2(_06744_ ), .ZN(_08338_ ) );
NAND3_X1 _23361_ ( .A1(_08247_ ), .A2(\u_lsu.pmem[2784] ), .A3(\alu_result_out[2] ), .ZN(_08339_ ) );
NAND4_X1 _23362_ ( .A1(_08337_ ), .A2(_08312_ ), .A3(_08338_ ), .A4(_08339_ ), .ZN(_08340_ ) );
NAND3_X1 _23363_ ( .A1(_09888_ ), .A2(_08335_ ), .A3(_08340_ ), .ZN(_08341_ ) );
NAND3_X1 _23364_ ( .A1(_08329_ ), .A2(_09785_ ), .A3(_08341_ ), .ZN(_08342_ ) );
AOI22_X1 _23365_ ( .A1(\u_lsu.pmem[2400] ), .A2(_08330_ ), .B1(_08242_ ), .B2(\u_lsu.pmem[2368] ), .ZN(_08343_ ) );
AOI22_X1 _23366_ ( .A1(\u_lsu.pmem[2336] ), .A2(_08331_ ), .B1(_09531_ ), .B2(\u_lsu.pmem[2304] ), .ZN(_08344_ ) );
NAND3_X1 _23367_ ( .A1(_08343_ ), .A2(_07009_ ), .A3(_08344_ ), .ZN(_08345_ ) );
AOI22_X1 _23368_ ( .A1(\u_lsu.pmem[2528] ), .A2(_08330_ ), .B1(_08242_ ), .B2(\u_lsu.pmem[2496] ), .ZN(_08346_ ) );
AOI22_X1 _23369_ ( .A1(\u_lsu.pmem[2464] ), .A2(_08331_ ), .B1(_09531_ ), .B2(\u_lsu.pmem[2432] ), .ZN(_08347_ ) );
NAND3_X1 _23370_ ( .A1(_08346_ ), .A2(\alu_result_out[4] ), .A3(_08347_ ), .ZN(_08348_ ) );
NAND3_X1 _23371_ ( .A1(\alu_result_out[5] ), .A2(_08345_ ), .A3(_08348_ ), .ZN(_08349_ ) );
AOI22_X1 _23372_ ( .A1(_08242_ ), .A2(\u_lsu.pmem[2112] ), .B1(_08336_ ), .B2(\u_lsu.pmem[2080] ), .ZN(_08350_ ) );
AOI22_X1 _23373_ ( .A1(_08251_ ), .A2(\u_lsu.pmem[2144] ), .B1(_08243_ ), .B2(\u_lsu.pmem[2048] ), .ZN(_08351_ ) );
AOI21_X1 _23374_ ( .A(_08231_ ), .B1(_08350_ ), .B2(_08351_ ), .ZN(_08352_ ) );
BUF_X4 _23375_ ( .A(_06339_ ), .Z(_08353_ ) );
AOI22_X1 _23376_ ( .A1(_08242_ ), .A2(\u_lsu.pmem[2240] ), .B1(_08353_ ), .B2(\u_lsu.pmem[2208] ), .ZN(_08354_ ) );
BUF_X4 _23377_ ( .A(_09530_ ), .Z(_08355_ ) );
AOI22_X1 _23378_ ( .A1(_08250_ ), .A2(\u_lsu.pmem[2272] ), .B1(_08355_ ), .B2(\u_lsu.pmem[2176] ), .ZN(_08356_ ) );
AOI21_X1 _23379_ ( .A(_07008_ ), .B1(_08354_ ), .B2(_08356_ ), .ZN(_08357_ ) );
OAI21_X1 _23380_ ( .A(_09888_ ), .B1(_08352_ ), .B2(_08357_ ), .ZN(_08358_ ) );
NAND3_X1 _23381_ ( .A1(_08349_ ), .A2(_09666_ ), .A3(_08358_ ), .ZN(_08359_ ) );
NAND3_X1 _23382_ ( .A1(_08342_ ), .A2(_09805_ ), .A3(_08359_ ), .ZN(_08360_ ) );
OAI211_X1 _23383_ ( .A(_06400_ ), .B(\u_lsu.pmem[4000] ), .C1(_06352_ ), .C2(_06355_ ), .ZN(_08361_ ) );
INV_X1 _23384_ ( .A(_08361_ ), .ZN(_08362_ ) );
AOI221_X4 _23385_ ( .A(_08362_ ), .B1(_06380_ ), .B2(\u_lsu.pmem[3968] ), .C1(\u_lsu.pmem[4064] ), .C2(_06316_ ), .ZN(_08363_ ) );
NAND3_X1 _23386_ ( .A1(\alu_result_out[3] ), .A2(_09096_ ), .A3(\u_lsu.pmem[4032] ), .ZN(_08364_ ) );
AOI21_X1 _23387_ ( .A(_08241_ ), .B1(_08363_ ), .B2(_08364_ ), .ZN(_08365_ ) );
OAI211_X1 _23388_ ( .A(_06436_ ), .B(\u_lsu.pmem[3872] ), .C1(_06351_ ), .C2(_06355_ ), .ZN(_08366_ ) );
INV_X1 _23389_ ( .A(_08366_ ), .ZN(_08367_ ) );
AOI221_X4 _23390_ ( .A(_08367_ ), .B1(_06221_ ), .B2(\u_lsu.pmem[3840] ), .C1(\u_lsu.pmem[3936] ), .C2(_06857_ ), .ZN(_08368_ ) );
NAND3_X1 _23391_ ( .A1(_08247_ ), .A2(_08283_ ), .A3(\u_lsu.pmem[3904] ), .ZN(_08369_ ) );
AOI21_X1 _23392_ ( .A(_08231_ ), .B1(_08368_ ), .B2(_08369_ ), .ZN(_08370_ ) );
OAI21_X1 _23393_ ( .A(\alu_result_out[5] ), .B1(_08365_ ), .B2(_08370_ ), .ZN(_08371_ ) );
AND3_X1 _23394_ ( .A1(_06434_ ), .A2(\u_lsu.pmem[3808] ), .A3(_06543_ ), .ZN(_08372_ ) );
AOI221_X4 _23395_ ( .A(_08372_ ), .B1(\u_lsu.pmem[3712] ), .B2(_06268_ ), .C1(\u_lsu.pmem[3776] ), .C2(_06469_ ), .ZN(_08373_ ) );
NAND3_X1 _23396_ ( .A1(_10433_ ), .A2(\u_lsu.pmem[3744] ), .A3(\alu_result_out[2] ), .ZN(_08374_ ) );
NAND3_X1 _23397_ ( .A1(_08373_ ), .A2(_08312_ ), .A3(_08374_ ), .ZN(_08375_ ) );
MUX2_X1 _23398_ ( .A(\u_lsu.pmem[3648] ), .B(\u_lsu.pmem[3680] ), .S(_06544_ ), .Z(_08376_ ) );
MUX2_X1 _23399_ ( .A(\u_lsu.pmem[3584] ), .B(\u_lsu.pmem[3616] ), .S(_06437_ ), .Z(_08377_ ) );
MUX2_X1 _23400_ ( .A(_08376_ ), .B(_08377_ ), .S(_10432_ ), .Z(_08378_ ) );
OAI211_X1 _23401_ ( .A(_08375_ ), .B(_08236_ ), .C1(\alu_result_out[4] ), .C2(_08378_ ), .ZN(_08379_ ) );
NAND3_X1 _23402_ ( .A1(_08371_ ), .A2(_08379_ ), .A3(_09785_ ), .ZN(_08380_ ) );
AOI22_X1 _23403_ ( .A1(\u_lsu.pmem[3424] ), .A2(_08330_ ), .B1(_08242_ ), .B2(\u_lsu.pmem[3392] ), .ZN(_08381_ ) );
AOI22_X1 _23404_ ( .A1(\u_lsu.pmem[3360] ), .A2(_08331_ ), .B1(_09531_ ), .B2(\u_lsu.pmem[3328] ), .ZN(_08382_ ) );
NAND3_X1 _23405_ ( .A1(_08381_ ), .A2(_07009_ ), .A3(_08382_ ), .ZN(_08383_ ) );
BUF_X4 _23406_ ( .A(_06741_ ), .Z(_08384_ ) );
AOI22_X1 _23407_ ( .A1(\u_lsu.pmem[3552] ), .A2(_08330_ ), .B1(_08384_ ), .B2(\u_lsu.pmem[3520] ), .ZN(_08385_ ) );
AOI22_X1 _23408_ ( .A1(\u_lsu.pmem[3488] ), .A2(_08331_ ), .B1(_09531_ ), .B2(\u_lsu.pmem[3456] ), .ZN(_08386_ ) );
NAND3_X1 _23409_ ( .A1(_08385_ ), .A2(\alu_result_out[4] ), .A3(_08386_ ), .ZN(_08387_ ) );
NAND3_X1 _23410_ ( .A1(\alu_result_out[5] ), .A2(_08383_ ), .A3(_08387_ ), .ZN(_08388_ ) );
AOI22_X1 _23411_ ( .A1(\u_lsu.pmem[3168] ), .A2(_08250_ ), .B1(_06741_ ), .B2(\u_lsu.pmem[3136] ), .ZN(_08389_ ) );
AOI22_X1 _23412_ ( .A1(\u_lsu.pmem[3104] ), .A2(_08336_ ), .B1(_08355_ ), .B2(\u_lsu.pmem[3072] ), .ZN(_08390_ ) );
AOI21_X1 _23413_ ( .A(_06721_ ), .B1(_08389_ ), .B2(_08390_ ), .ZN(_08391_ ) );
AOI22_X1 _23414_ ( .A1(\u_lsu.pmem[3296] ), .A2(_08250_ ), .B1(_06741_ ), .B2(\u_lsu.pmem[3264] ), .ZN(_08392_ ) );
AOI22_X1 _23415_ ( .A1(\u_lsu.pmem[3232] ), .A2(_08353_ ), .B1(_09530_ ), .B2(\u_lsu.pmem[3200] ), .ZN(_08393_ ) );
AOI21_X1 _23416_ ( .A(_07008_ ), .B1(_08392_ ), .B2(_08393_ ), .ZN(_08394_ ) );
OAI21_X1 _23417_ ( .A(_08236_ ), .B1(_08391_ ), .B2(_08394_ ), .ZN(_08395_ ) );
NAND3_X1 _23418_ ( .A1(_08388_ ), .A2(_09666_ ), .A3(_08395_ ), .ZN(_08396_ ) );
NAND3_X1 _23419_ ( .A1(_08380_ ), .A2(_10286_ ), .A3(_08396_ ), .ZN(_08397_ ) );
NAND3_X1 _23420_ ( .A1(_08360_ ), .A2(_09605_ ), .A3(_08397_ ), .ZN(_08398_ ) );
NAND3_X1 _23421_ ( .A1(_08321_ ), .A2(_02481_ ), .A3(_08398_ ), .ZN(_08399_ ) );
AND3_X1 _23422_ ( .A1(_06440_ ), .A2(\u_lsu.pmem[7712] ), .A3(_06436_ ), .ZN(_08400_ ) );
AOI221_X4 _23423_ ( .A(_08400_ ), .B1(\u_lsu.pmem[7680] ), .B2(_06524_ ), .C1(\u_lsu.pmem[7776] ), .C2(_06605_ ), .ZN(_08401_ ) );
NAND3_X1 _23424_ ( .A1(\alu_result_out[3] ), .A2(_09096_ ), .A3(\u_lsu.pmem[7744] ), .ZN(_08402_ ) );
AOI21_X1 _23425_ ( .A(_08312_ ), .B1(_08401_ ), .B2(_08402_ ), .ZN(_08403_ ) );
AND3_X1 _23426_ ( .A1(_10430_ ), .A2(\u_lsu.pmem[7840] ), .A3(_06543_ ), .ZN(_08404_ ) );
AOI221_X4 _23427_ ( .A(_08404_ ), .B1(\u_lsu.pmem[7808] ), .B2(_06445_ ), .C1(\u_lsu.pmem[7904] ), .C2(_06637_ ), .ZN(_08405_ ) );
NAND3_X1 _23428_ ( .A1(_08247_ ), .A2(_08283_ ), .A3(\u_lsu.pmem[7872] ), .ZN(_08406_ ) );
AOI21_X1 _23429_ ( .A(_07008_ ), .B1(_08405_ ), .B2(_08406_ ), .ZN(_08407_ ) );
OAI21_X1 _23430_ ( .A(_09888_ ), .B1(_08403_ ), .B2(_08407_ ), .ZN(_08408_ ) );
AOI22_X1 _23431_ ( .A1(_06593_ ), .A2(\u_lsu.pmem[8128] ), .B1(_06794_ ), .B2(\u_lsu.pmem[8096] ), .ZN(_08409_ ) );
NAND3_X1 _23432_ ( .A1(_06619_ ), .A2(\u_lsu.pmem[8160] ), .A3(_06249_ ), .ZN(_08410_ ) );
OAI211_X1 _23433_ ( .A(_06515_ ), .B(\u_lsu.pmem[8064] ), .C1(_06587_ ), .C2(_06588_ ), .ZN(_08411_ ) );
AND4_X1 _23434_ ( .A1(_06234_ ), .A2(_08409_ ), .A3(_08410_ ), .A4(_08411_ ), .ZN(_08412_ ) );
AOI22_X1 _23435_ ( .A1(_06836_ ), .A2(\u_lsu.pmem[8000] ), .B1(_06640_ ), .B2(\u_lsu.pmem[7936] ), .ZN(_08413_ ) );
NAND3_X1 _23436_ ( .A1(_06473_ ), .A2(\u_lsu.pmem[8032] ), .A3(_06333_ ), .ZN(_08414_ ) );
OAI211_X1 _23437_ ( .A(_06401_ ), .B(\u_lsu.pmem[7968] ), .C1(_06480_ ), .C2(_06481_ ), .ZN(_08415_ ) );
AND4_X1 _23438_ ( .A1(_06479_ ), .A2(_08413_ ), .A3(_08414_ ), .A4(_08415_ ), .ZN(_08416_ ) );
OR3_X1 _23439_ ( .A1(_08412_ ), .A2(_08416_ ), .A3(_09744_ ), .ZN(_08417_ ) );
AOI21_X1 _23440_ ( .A(_09666_ ), .B1(_08408_ ), .B2(_08417_ ), .ZN(_08418_ ) );
AOI22_X1 _23441_ ( .A1(\u_lsu.pmem[7520] ), .A2(_08330_ ), .B1(_08384_ ), .B2(\u_lsu.pmem[7488] ), .ZN(_08419_ ) );
AOI22_X1 _23442_ ( .A1(\u_lsu.pmem[7456] ), .A2(_08336_ ), .B1(_08243_ ), .B2(\u_lsu.pmem[7424] ), .ZN(_08420_ ) );
NAND3_X1 _23443_ ( .A1(_08419_ ), .A2(_08241_ ), .A3(_08420_ ), .ZN(_08421_ ) );
AOI22_X1 _23444_ ( .A1(\u_lsu.pmem[7648] ), .A2(_08251_ ), .B1(_06741_ ), .B2(\u_lsu.pmem[7616] ), .ZN(_08422_ ) );
AOI22_X1 _23445_ ( .A1(\u_lsu.pmem[7584] ), .A2(_08336_ ), .B1(_08243_ ), .B2(\u_lsu.pmem[7552] ), .ZN(_08423_ ) );
NAND3_X1 _23446_ ( .A1(_08422_ ), .A2(_08312_ ), .A3(_08423_ ), .ZN(_08424_ ) );
NAND3_X1 _23447_ ( .A1(_10529_ ), .A2(_08421_ ), .A3(_08424_ ), .ZN(_08425_ ) );
AOI22_X1 _23448_ ( .A1(\u_lsu.pmem[7264] ), .A2(_08251_ ), .B1(_06741_ ), .B2(\u_lsu.pmem[7232] ), .ZN(_08426_ ) );
AOI22_X1 _23449_ ( .A1(\u_lsu.pmem[7200] ), .A2(_08336_ ), .B1(_08355_ ), .B2(\u_lsu.pmem[7168] ), .ZN(_08427_ ) );
NAND3_X1 _23450_ ( .A1(_08426_ ), .A2(_08241_ ), .A3(_08427_ ), .ZN(_08428_ ) );
AOI22_X1 _23451_ ( .A1(\u_lsu.pmem[7392] ), .A2(_08251_ ), .B1(_06741_ ), .B2(\u_lsu.pmem[7360] ), .ZN(_08429_ ) );
AOI22_X1 _23452_ ( .A1(\u_lsu.pmem[7328] ), .A2(_08353_ ), .B1(_08355_ ), .B2(\u_lsu.pmem[7296] ), .ZN(_08430_ ) );
NAND3_X1 _23453_ ( .A1(_08429_ ), .A2(_08312_ ), .A3(_08430_ ), .ZN(_08431_ ) );
NAND3_X1 _23454_ ( .A1(_08236_ ), .A2(_08428_ ), .A3(_08431_ ), .ZN(_08432_ ) );
AOI21_X1 _23455_ ( .A(_09784_ ), .B1(_08425_ ), .B2(_08432_ ), .ZN(_08433_ ) );
OAI21_X1 _23456_ ( .A(_10286_ ), .B1(_08418_ ), .B2(_08433_ ), .ZN(_08434_ ) );
AND3_X1 _23457_ ( .A1(_06434_ ), .A2(_06598_ ), .A3(\u_lsu.pmem[6336] ), .ZN(_08435_ ) );
AOI221_X4 _23458_ ( .A(_08435_ ), .B1(\u_lsu.pmem[6304] ), .B2(_06264_ ), .C1(\u_lsu.pmem[6272] ), .C2(_09530_ ), .ZN(_08436_ ) );
NAND3_X1 _23459_ ( .A1(\alu_result_out[3] ), .A2(\u_lsu.pmem[6368] ), .A3(\alu_result_out[2] ), .ZN(_08437_ ) );
NAND3_X1 _23460_ ( .A1(_08436_ ), .A2(_08312_ ), .A3(_08437_ ), .ZN(_08438_ ) );
MUX2_X1 _23461_ ( .A(\u_lsu.pmem[6208] ), .B(\u_lsu.pmem[6240] ), .S(_06408_ ), .Z(_08439_ ) );
MUX2_X1 _23462_ ( .A(\u_lsu.pmem[6144] ), .B(\u_lsu.pmem[6176] ), .S(_06408_ ), .Z(_08440_ ) );
MUX2_X1 _23463_ ( .A(_08439_ ), .B(_08440_ ), .S(_10432_ ), .Z(_08441_ ) );
OAI211_X1 _23464_ ( .A(_08438_ ), .B(_08236_ ), .C1(\alu_result_out[4] ), .C2(_08441_ ), .ZN(_08442_ ) );
AOI22_X1 _23465_ ( .A1(\u_lsu.pmem[6624] ), .A2(_08251_ ), .B1(_08384_ ), .B2(\u_lsu.pmem[6592] ), .ZN(_08443_ ) );
AOI22_X1 _23466_ ( .A1(\u_lsu.pmem[6560] ), .A2(_08331_ ), .B1(_09531_ ), .B2(\u_lsu.pmem[6528] ), .ZN(_08444_ ) );
AOI21_X1 _23467_ ( .A(_08241_ ), .B1(_08443_ ), .B2(_08444_ ), .ZN(_08445_ ) );
AOI22_X1 _23468_ ( .A1(\u_lsu.pmem[6496] ), .A2(_08250_ ), .B1(_06741_ ), .B2(\u_lsu.pmem[6464] ), .ZN(_08446_ ) );
AOI22_X1 _23469_ ( .A1(\u_lsu.pmem[6432] ), .A2(_08336_ ), .B1(_08355_ ), .B2(\u_lsu.pmem[6400] ), .ZN(_08447_ ) );
AOI21_X1 _23470_ ( .A(_06721_ ), .B1(_08446_ ), .B2(_08447_ ), .ZN(_08448_ ) );
OAI21_X1 _23471_ ( .A(_10529_ ), .B1(_08445_ ), .B2(_08448_ ), .ZN(_08449_ ) );
NAND3_X1 _23472_ ( .A1(_08442_ ), .A2(_09666_ ), .A3(_08449_ ), .ZN(_08450_ ) );
OAI211_X1 _23473_ ( .A(_06400_ ), .B(\u_lsu.pmem[6944] ), .C1(_06352_ ), .C2(_06355_ ), .ZN(_08451_ ) );
INV_X1 _23474_ ( .A(_08451_ ), .ZN(_08452_ ) );
AOI221_X4 _23475_ ( .A(_08452_ ), .B1(_06274_ ), .B2(\u_lsu.pmem[6912] ), .C1(\u_lsu.pmem[7008] ), .C2(_06605_ ), .ZN(_08453_ ) );
NAND3_X1 _23476_ ( .A1(\alu_result_out[3] ), .A2(_09096_ ), .A3(\u_lsu.pmem[6976] ), .ZN(_08454_ ) );
AOI21_X1 _23477_ ( .A(_08312_ ), .B1(_08453_ ), .B2(_08454_ ), .ZN(_08455_ ) );
AOI22_X1 _23478_ ( .A1(_08242_ ), .A2(\u_lsu.pmem[7104] ), .B1(_08353_ ), .B2(\u_lsu.pmem[7072] ), .ZN(_08456_ ) );
AOI22_X1 _23479_ ( .A1(_08251_ ), .A2(\u_lsu.pmem[7136] ), .B1(_08355_ ), .B2(\u_lsu.pmem[7040] ), .ZN(_08457_ ) );
AOI21_X1 _23480_ ( .A(_07008_ ), .B1(_08456_ ), .B2(_08457_ ), .ZN(_08458_ ) );
OAI21_X1 _23481_ ( .A(\alu_result_out[5] ), .B1(_08455_ ), .B2(_08458_ ), .ZN(_08459_ ) );
AOI22_X1 _23482_ ( .A1(\u_lsu.pmem[6752] ), .A2(_08330_ ), .B1(_08384_ ), .B2(\u_lsu.pmem[6720] ), .ZN(_08460_ ) );
AOI22_X1 _23483_ ( .A1(\u_lsu.pmem[6688] ), .A2(_08331_ ), .B1(_09531_ ), .B2(\u_lsu.pmem[6656] ), .ZN(_08461_ ) );
NAND3_X1 _23484_ ( .A1(_08460_ ), .A2(_07009_ ), .A3(_08461_ ), .ZN(_08462_ ) );
AOI22_X1 _23485_ ( .A1(\u_lsu.pmem[6880] ), .A2(_08330_ ), .B1(_08384_ ), .B2(\u_lsu.pmem[6848] ), .ZN(_08463_ ) );
AOI22_X1 _23486_ ( .A1(\u_lsu.pmem[6816] ), .A2(_08336_ ), .B1(_08243_ ), .B2(\u_lsu.pmem[6784] ), .ZN(_08464_ ) );
NAND3_X1 _23487_ ( .A1(_08463_ ), .A2(_08312_ ), .A3(_08464_ ), .ZN(_08465_ ) );
NAND3_X1 _23488_ ( .A1(_09888_ ), .A2(_08462_ ), .A3(_08465_ ), .ZN(_08466_ ) );
NAND3_X1 _23489_ ( .A1(_08459_ ), .A2(_09785_ ), .A3(_08466_ ), .ZN(_08467_ ) );
NAND3_X1 _23490_ ( .A1(_08450_ ), .A2(_08467_ ), .A3(_09805_ ), .ZN(_08468_ ) );
NAND3_X1 _23491_ ( .A1(_08434_ ), .A2(_09605_ ), .A3(_08468_ ), .ZN(_08469_ ) );
AOI22_X1 _23492_ ( .A1(_08251_ ), .A2(\u_lsu.pmem[5088] ), .B1(_08353_ ), .B2(\u_lsu.pmem[5024] ), .ZN(_08470_ ) );
NAND3_X1 _23493_ ( .A1(_10433_ ), .A2(\u_lsu.pmem[4992] ), .A3(_08283_ ), .ZN(_08471_ ) );
NAND3_X1 _23494_ ( .A1(_08232_ ), .A2(_08233_ ), .A3(\u_lsu.pmem[5056] ), .ZN(_08472_ ) );
NAND4_X1 _23495_ ( .A1(_08470_ ), .A2(_08231_ ), .A3(_08471_ ), .A4(_08472_ ), .ZN(_08473_ ) );
AOI22_X1 _23496_ ( .A1(_08242_ ), .A2(\u_lsu.pmem[4928] ), .B1(_08243_ ), .B2(\u_lsu.pmem[4864] ), .ZN(_08474_ ) );
NAND3_X1 _23497_ ( .A1(_08232_ ), .A2(\u_lsu.pmem[4960] ), .A3(\alu_result_out[2] ), .ZN(_08475_ ) );
NAND3_X1 _23498_ ( .A1(_10433_ ), .A2(\u_lsu.pmem[4896] ), .A3(_08245_ ), .ZN(_08476_ ) );
NAND4_X1 _23499_ ( .A1(_08474_ ), .A2(_08241_ ), .A3(_08475_ ), .A4(_08476_ ), .ZN(_08477_ ) );
NAND3_X1 _23500_ ( .A1(_10529_ ), .A2(_08473_ ), .A3(_08477_ ), .ZN(_08478_ ) );
AOI22_X1 _23501_ ( .A1(_08251_ ), .A2(\u_lsu.pmem[4704] ), .B1(_08355_ ), .B2(\u_lsu.pmem[4608] ), .ZN(_08479_ ) );
OAI211_X1 _23502_ ( .A(_06675_ ), .B(\u_lsu.pmem[4640] ), .C1(_06743_ ), .C2(_06744_ ), .ZN(_08480_ ) );
NAND3_X1 _23503_ ( .A1(_08232_ ), .A2(_08233_ ), .A3(\u_lsu.pmem[4672] ), .ZN(_08481_ ) );
NAND4_X1 _23504_ ( .A1(_08479_ ), .A2(_08241_ ), .A3(_08480_ ), .A4(_08481_ ), .ZN(_08482_ ) );
AOI22_X1 _23505_ ( .A1(_08250_ ), .A2(\u_lsu.pmem[4832] ), .B1(_08355_ ), .B2(\u_lsu.pmem[4736] ), .ZN(_08483_ ) );
OAI211_X1 _23506_ ( .A(_06675_ ), .B(\u_lsu.pmem[4768] ), .C1(_06743_ ), .C2(_06744_ ), .ZN(_08484_ ) );
NAND3_X1 _23507_ ( .A1(_08232_ ), .A2(_08233_ ), .A3(\u_lsu.pmem[4800] ), .ZN(_08485_ ) );
NAND4_X1 _23508_ ( .A1(_08483_ ), .A2(_08231_ ), .A3(_08484_ ), .A4(_08485_ ), .ZN(_08486_ ) );
NAND3_X1 _23509_ ( .A1(_08236_ ), .A2(_08482_ ), .A3(_08486_ ), .ZN(_08487_ ) );
AOI21_X1 _23510_ ( .A(_09666_ ), .B1(_08478_ ), .B2(_08487_ ), .ZN(_08488_ ) );
AOI22_X1 _23511_ ( .A1(_08384_ ), .A2(\u_lsu.pmem[4416] ), .B1(_08353_ ), .B2(\u_lsu.pmem[4384] ), .ZN(_08489_ ) );
OAI211_X1 _23512_ ( .A(_08233_ ), .B(\u_lsu.pmem[4352] ), .C1(_06743_ ), .C2(_06744_ ), .ZN(_08490_ ) );
NAND3_X1 _23513_ ( .A1(_09071_ ), .A2(\u_lsu.pmem[4448] ), .A3(_08245_ ), .ZN(_08491_ ) );
NAND4_X1 _23514_ ( .A1(_08489_ ), .A2(_07008_ ), .A3(_08490_ ), .A4(_08491_ ), .ZN(_08492_ ) );
AOI22_X1 _23515_ ( .A1(_08384_ ), .A2(\u_lsu.pmem[4544] ), .B1(_08353_ ), .B2(\u_lsu.pmem[4512] ), .ZN(_08493_ ) );
OAI211_X1 _23516_ ( .A(_08233_ ), .B(\u_lsu.pmem[4480] ), .C1(_06743_ ), .C2(_06744_ ), .ZN(_08494_ ) );
NAND3_X1 _23517_ ( .A1(_09071_ ), .A2(\u_lsu.pmem[4576] ), .A3(_08245_ ), .ZN(_08495_ ) );
NAND4_X1 _23518_ ( .A1(_08493_ ), .A2(_06721_ ), .A3(_08494_ ), .A4(_08495_ ), .ZN(_08496_ ) );
NAND3_X1 _23519_ ( .A1(_10529_ ), .A2(_08492_ ), .A3(_08496_ ), .ZN(_08497_ ) );
AOI22_X1 _23520_ ( .A1(\u_lsu.pmem[4192] ), .A2(_08250_ ), .B1(_06741_ ), .B2(\u_lsu.pmem[4160] ), .ZN(_08498_ ) );
AOI22_X1 _23521_ ( .A1(\u_lsu.pmem[4128] ), .A2(_08353_ ), .B1(_08355_ ), .B2(\u_lsu.pmem[4096] ), .ZN(_08499_ ) );
NAND3_X1 _23522_ ( .A1(_08498_ ), .A2(_08241_ ), .A3(_08499_ ), .ZN(_08500_ ) );
AOI22_X1 _23523_ ( .A1(\u_lsu.pmem[4256] ), .A2(_08353_ ), .B1(_09530_ ), .B2(\u_lsu.pmem[4224] ), .ZN(_08501_ ) );
NAND3_X1 _23524_ ( .A1(_09071_ ), .A2(_08233_ ), .A3(\u_lsu.pmem[4288] ), .ZN(_08502_ ) );
NAND3_X1 _23525_ ( .A1(_09071_ ), .A2(\u_lsu.pmem[4320] ), .A3(_06675_ ), .ZN(_08503_ ) );
NAND4_X1 _23526_ ( .A1(_08501_ ), .A2(_06721_ ), .A3(_08502_ ), .A4(_08503_ ), .ZN(_08504_ ) );
NAND3_X1 _23527_ ( .A1(_08236_ ), .A2(_08500_ ), .A3(_08504_ ), .ZN(_08505_ ) );
AOI21_X1 _23528_ ( .A(_09784_ ), .B1(_08497_ ), .B2(_08505_ ), .ZN(_08506_ ) );
OAI21_X1 _23529_ ( .A(_09805_ ), .B1(_08488_ ), .B2(_08506_ ), .ZN(_08507_ ) );
AOI22_X1 _23530_ ( .A1(\u_lsu.pmem[5472] ), .A2(_08330_ ), .B1(_08242_ ), .B2(\u_lsu.pmem[5440] ), .ZN(_08508_ ) );
AOI22_X1 _23531_ ( .A1(\u_lsu.pmem[5408] ), .A2(_08331_ ), .B1(_09531_ ), .B2(\u_lsu.pmem[5376] ), .ZN(_08509_ ) );
NAND3_X1 _23532_ ( .A1(_08508_ ), .A2(_07009_ ), .A3(_08509_ ), .ZN(_08510_ ) );
AOI22_X1 _23533_ ( .A1(\u_lsu.pmem[5536] ), .A2(_08331_ ), .B1(_09531_ ), .B2(\u_lsu.pmem[5504] ), .ZN(_08511_ ) );
NAND3_X1 _23534_ ( .A1(_08247_ ), .A2(\u_lsu.pmem[5600] ), .A3(\alu_result_out[2] ), .ZN(_08512_ ) );
NAND3_X1 _23535_ ( .A1(_08247_ ), .A2(_08283_ ), .A3(\u_lsu.pmem[5568] ), .ZN(_08513_ ) );
NAND4_X1 _23536_ ( .A1(_08511_ ), .A2(_08312_ ), .A3(_08512_ ), .A4(_08513_ ), .ZN(_08514_ ) );
NAND3_X1 _23537_ ( .A1(\alu_result_out[5] ), .A2(_08510_ ), .A3(_08514_ ), .ZN(_08515_ ) );
AOI22_X1 _23538_ ( .A1(\u_lsu.pmem[5216] ), .A2(_08330_ ), .B1(_08384_ ), .B2(\u_lsu.pmem[5184] ), .ZN(_08516_ ) );
AOI22_X1 _23539_ ( .A1(\u_lsu.pmem[5152] ), .A2(_08336_ ), .B1(_08243_ ), .B2(\u_lsu.pmem[5120] ), .ZN(_08517_ ) );
NAND3_X1 _23540_ ( .A1(_08516_ ), .A2(_08241_ ), .A3(_08517_ ), .ZN(_08518_ ) );
AOI22_X1 _23541_ ( .A1(\u_lsu.pmem[5280] ), .A2(_08336_ ), .B1(_08243_ ), .B2(\u_lsu.pmem[5248] ), .ZN(_08519_ ) );
NAND3_X1 _23542_ ( .A1(_08232_ ), .A2(_08233_ ), .A3(\u_lsu.pmem[5312] ), .ZN(_08520_ ) );
NAND3_X1 _23543_ ( .A1(_08232_ ), .A2(\u_lsu.pmem[5344] ), .A3(_08245_ ), .ZN(_08521_ ) );
NAND4_X1 _23544_ ( .A1(_08519_ ), .A2(_08231_ ), .A3(_08520_ ), .A4(_08521_ ), .ZN(_08522_ ) );
NAND3_X1 _23545_ ( .A1(_08236_ ), .A2(_08518_ ), .A3(_08522_ ), .ZN(_08523_ ) );
NAND3_X1 _23546_ ( .A1(_08515_ ), .A2(_09666_ ), .A3(_08523_ ), .ZN(_08524_ ) );
AOI22_X1 _23547_ ( .A1(\u_lsu.pmem[5920] ), .A2(_08331_ ), .B1(_09531_ ), .B2(\u_lsu.pmem[5888] ), .ZN(_08525_ ) );
NAND3_X1 _23548_ ( .A1(_08247_ ), .A2(_08283_ ), .A3(\u_lsu.pmem[5952] ), .ZN(_08526_ ) );
NAND3_X1 _23549_ ( .A1(_08232_ ), .A2(\u_lsu.pmem[5984] ), .A3(\alu_result_out[2] ), .ZN(_08527_ ) );
NAND4_X1 _23550_ ( .A1(_08525_ ), .A2(_08241_ ), .A3(_08526_ ), .A4(_08527_ ), .ZN(_08528_ ) );
AOI22_X1 _23551_ ( .A1(_08251_ ), .A2(\u_lsu.pmem[6112] ), .B1(_08243_ ), .B2(\u_lsu.pmem[6016] ), .ZN(_08529_ ) );
NAND3_X1 _23552_ ( .A1(_08247_ ), .A2(_08283_ ), .A3(\u_lsu.pmem[6080] ), .ZN(_08530_ ) );
OAI211_X1 _23553_ ( .A(_08245_ ), .B(\u_lsu.pmem[6048] ), .C1(_06743_ ), .C2(_06744_ ), .ZN(_08531_ ) );
NAND4_X1 _23554_ ( .A1(_08529_ ), .A2(_08231_ ), .A3(_08530_ ), .A4(_08531_ ), .ZN(_08532_ ) );
NAND3_X1 _23555_ ( .A1(\alu_result_out[5] ), .A2(_08528_ ), .A3(_08532_ ), .ZN(_08533_ ) );
AOI22_X1 _23556_ ( .A1(_08384_ ), .A2(\u_lsu.pmem[5696] ), .B1(_08353_ ), .B2(\u_lsu.pmem[5664] ), .ZN(_08534_ ) );
NAND3_X1 _23557_ ( .A1(_08232_ ), .A2(\u_lsu.pmem[5728] ), .A3(_08245_ ), .ZN(_08535_ ) );
NAND3_X1 _23558_ ( .A1(_10433_ ), .A2(\u_lsu.pmem[5632] ), .A3(_08233_ ), .ZN(_08536_ ) );
NAND4_X1 _23559_ ( .A1(_08534_ ), .A2(_07008_ ), .A3(_08535_ ), .A4(_08536_ ), .ZN(_08537_ ) );
AOI22_X1 _23560_ ( .A1(_08384_ ), .A2(\u_lsu.pmem[5824] ), .B1(_08355_ ), .B2(\u_lsu.pmem[5760] ), .ZN(_08538_ ) );
NAND3_X1 _23561_ ( .A1(_10433_ ), .A2(\u_lsu.pmem[5792] ), .A3(_08245_ ), .ZN(_08539_ ) );
NAND3_X1 _23562_ ( .A1(_09071_ ), .A2(\u_lsu.pmem[5856] ), .A3(_08245_ ), .ZN(_08540_ ) );
NAND4_X1 _23563_ ( .A1(_08538_ ), .A2(_08231_ ), .A3(_08539_ ), .A4(_08540_ ), .ZN(_08541_ ) );
NAND3_X1 _23564_ ( .A1(_08236_ ), .A2(_08537_ ), .A3(_08541_ ), .ZN(_08542_ ) );
NAND3_X1 _23565_ ( .A1(_08533_ ), .A2(_09785_ ), .A3(_08542_ ), .ZN(_08543_ ) );
NAND3_X1 _23566_ ( .A1(_08524_ ), .A2(_08543_ ), .A3(_10286_ ), .ZN(_08544_ ) );
NAND3_X1 _23567_ ( .A1(_08507_ ), .A2(_02484_ ), .A3(_08544_ ), .ZN(_08545_ ) );
NAND3_X1 _23568_ ( .A1(_08469_ ), .A2(_10045_ ), .A3(_08545_ ), .ZN(_08546_ ) );
AOI21_X1 _23569_ ( .A(_05735_ ), .B1(_08399_ ), .B2(_08546_ ), .ZN(\load_data_out[0] ) );
XOR2_X1 _23570_ ( .A(_08954_ ), .B(_08955_ ), .Z(\alu_result_out[0] ) );
AND3_X1 _23571_ ( .A1(\alu_result_out[0] ), .A2(_06078_ ), .A3(_05735_ ), .ZN(_08547_ ) );
OAI21_X1 _23572_ ( .A(_06102_ ), .B1(\load_data_out[0] ), .B2(_08547_ ), .ZN(_08548_ ) );
AOI22_X1 _23573_ ( .A1(\alu_result_out[0] ), .A2(_06081_ ), .B1(\pc_out[0] ), .B2(_08908_ ), .ZN(_08549_ ) );
AOI21_X1 _23574_ ( .A(_06076_ ), .B1(_08548_ ), .B2(_08549_ ), .ZN(_00030_ ) );
AND2_X1 _23575_ ( .A1(\alu_result_out[27] ), .A2(_06078_ ), .ZN(_08550_ ) );
OAI21_X1 _23576_ ( .A(_06065_ ), .B1(_06077_ ), .B2(_08550_ ), .ZN(_08551_ ) );
NAND2_X1 _23577_ ( .A1(\alu_result_out[27] ), .A2(_06081_ ), .ZN(_08552_ ) );
OR2_X1 _23578_ ( .A1(_09391_ ), .A2(_08928_ ), .ZN(_08553_ ) );
AND3_X2 _23579_ ( .A1(_08551_ ), .A2(_08552_ ), .A3(_08553_ ), .ZN(_08554_ ) );
NOR2_X1 _23580_ ( .A1(_08554_ ), .A2(_06137_ ), .ZN(_00031_ ) );
AOI22_X1 _23581_ ( .A1(\alu_result_out[26] ), .A2(_06088_ ), .B1(_06082_ ), .B2(_09394_ ), .ZN(_08555_ ) );
AOI21_X1 _23582_ ( .A(_06076_ ), .B1(_06092_ ), .B2(_08555_ ), .ZN(_00032_ ) );
AOI22_X1 _23583_ ( .A1(\alu_result_out[25] ), .A2(_06088_ ), .B1(_06082_ ), .B2(_09403_ ), .ZN(_08556_ ) );
AOI21_X1 _23584_ ( .A(_06074_ ), .B1(_06092_ ), .B2(_08556_ ), .ZN(_00033_ ) );
AOI22_X1 _23585_ ( .A1(\alu_result_out[24] ), .A2(_06088_ ), .B1(_08908_ ), .B2(_09407_ ), .ZN(_08557_ ) );
AOI21_X1 _23586_ ( .A(_06074_ ), .B1(_06092_ ), .B2(_08557_ ), .ZN(_00034_ ) );
AND2_X1 _23587_ ( .A1(\alu_result_out[23] ), .A2(_06078_ ), .ZN(_08558_ ) );
OAI21_X1 _23588_ ( .A(_06065_ ), .B1(_06077_ ), .B2(_08558_ ), .ZN(_08559_ ) );
NAND2_X1 _23589_ ( .A1(\alu_result_out[23] ), .A2(_06081_ ), .ZN(_08560_ ) );
OR2_X1 _23590_ ( .A1(_09417_ ), .A2(_08928_ ), .ZN(_08561_ ) );
AND3_X2 _23591_ ( .A1(_08559_ ), .A2(_08560_ ), .A3(_08561_ ), .ZN(_08562_ ) );
NOR2_X1 _23592_ ( .A1(_08562_ ), .A2(_06137_ ), .ZN(_00035_ ) );
AOI22_X1 _23593_ ( .A1(\alu_result_out[22] ), .A2(_06088_ ), .B1(_08908_ ), .B2(_09419_ ), .ZN(_08563_ ) );
AOI21_X1 _23594_ ( .A(_06074_ ), .B1(_06092_ ), .B2(_08563_ ), .ZN(_00036_ ) );
NOR2_X1 _23595_ ( .A1(_06070_ ), .A2(\ifu_rdata[7] ), .ZN(_08564_ ) );
NAND2_X2 _23596_ ( .A1(_06072_ ), .A2(_08564_ ), .ZN(_08565_ ) );
BUF_X4 _23597_ ( .A(_08565_ ), .Z(_08566_ ) );
NOR2_X1 _23598_ ( .A1(_06066_ ), .A2(_08566_ ), .ZN(_00037_ ) );
BUF_X4 _23599_ ( .A(_08565_ ), .Z(_08567_ ) );
AOI21_X1 _23600_ ( .A(_08567_ ), .B1(_06080_ ), .B2(_06083_ ), .ZN(_00038_ ) );
NOR2_X1 _23601_ ( .A1(_06090_ ), .A2(_08566_ ), .ZN(_00039_ ) );
AOI21_X1 _23602_ ( .A(_08567_ ), .B1(_06092_ ), .B2(_06093_ ), .ZN(_00040_ ) );
NOR2_X1 _23603_ ( .A1(_06096_ ), .A2(_08566_ ), .ZN(_00041_ ) );
AOI21_X1 _23604_ ( .A(_08567_ ), .B1(_06092_ ), .B2(_06097_ ), .ZN(_00042_ ) );
NOR2_X1 _23605_ ( .A1(_06100_ ), .A2(_08566_ ), .ZN(_00043_ ) );
AOI21_X1 _23606_ ( .A(_08567_ ), .B1(_06104_ ), .B2(_06105_ ), .ZN(_00044_ ) );
NOR2_X1 _23607_ ( .A1(_06110_ ), .A2(_08566_ ), .ZN(_00045_ ) );
BUF_X4 _23608_ ( .A(_06091_ ), .Z(_08568_ ) );
AOI21_X1 _23609_ ( .A(_08567_ ), .B1(_08568_ ), .B2(_06111_ ), .ZN(_00046_ ) );
AOI21_X1 _23610_ ( .A(_08567_ ), .B1(_08568_ ), .B2(_06112_ ), .ZN(_00047_ ) );
AOI21_X1 _23611_ ( .A(_08567_ ), .B1(_06114_ ), .B2(_06115_ ), .ZN(_00048_ ) );
NOR2_X1 _23612_ ( .A1(_06120_ ), .A2(_08566_ ), .ZN(_00049_ ) );
NOR2_X1 _23613_ ( .A1(_06123_ ), .A2(_08566_ ), .ZN(_00050_ ) );
NOR2_X1 _23614_ ( .A1(_06128_ ), .A2(_08566_ ), .ZN(_00051_ ) );
NOR2_X1 _23615_ ( .A1(_06132_ ), .A2(_08566_ ), .ZN(_00052_ ) );
BUF_X4 _23616_ ( .A(_08565_ ), .Z(_08569_ ) );
NOR2_X1 _23617_ ( .A1(_06136_ ), .A2(_08569_ ), .ZN(_00053_ ) );
NOR2_X1 _23618_ ( .A1(_06140_ ), .A2(_08569_ ), .ZN(_00054_ ) );
NOR2_X1 _23619_ ( .A1(_06669_ ), .A2(_08569_ ), .ZN(_00055_ ) );
NOR2_X1 _23620_ ( .A1(_07007_ ), .A2(_08569_ ), .ZN(_00056_ ) );
NOR2_X1 _23621_ ( .A1(_07315_ ), .A2(_08569_ ), .ZN(_00057_ ) );
NOR2_X1 _23622_ ( .A1(_07617_ ), .A2(_08569_ ), .ZN(_00058_ ) );
NOR2_X1 _23623_ ( .A1(_07913_ ), .A2(_08569_ ), .ZN(_00059_ ) );
AOI21_X1 _23624_ ( .A(_08567_ ), .B1(_07915_ ), .B2(_07916_ ), .ZN(_00060_ ) );
NOR2_X1 _23625_ ( .A1(_08228_ ), .A2(_08569_ ), .ZN(_00061_ ) );
AOI21_X1 _23626_ ( .A(_08567_ ), .B1(_08548_ ), .B2(_08549_ ), .ZN(_00062_ ) );
NOR2_X1 _23627_ ( .A1(_08554_ ), .A2(_08569_ ), .ZN(_00063_ ) );
AOI21_X1 _23628_ ( .A(_08567_ ), .B1(_08568_ ), .B2(_08555_ ), .ZN(_00064_ ) );
AOI21_X1 _23629_ ( .A(_08565_ ), .B1(_08568_ ), .B2(_08556_ ), .ZN(_00065_ ) );
AOI21_X1 _23630_ ( .A(_08565_ ), .B1(_08568_ ), .B2(_08557_ ), .ZN(_00066_ ) );
NOR2_X1 _23631_ ( .A1(_08562_ ), .A2(_08569_ ), .ZN(_00067_ ) );
AOI21_X1 _23632_ ( .A(_08565_ ), .B1(_08568_ ), .B2(_08563_ ), .ZN(_00068_ ) );
AND3_X1 _23633_ ( .A1(_08586_ ), .A2(\ifu_rdata[7] ), .A3(\ifu_rdata[8] ), .ZN(_08570_ ) );
NAND2_X2 _23634_ ( .A1(_06068_ ), .A2(_08570_ ), .ZN(_08571_ ) );
BUF_X4 _23635_ ( .A(_08571_ ), .Z(_08572_ ) );
NOR2_X1 _23636_ ( .A1(_06066_ ), .A2(_08572_ ), .ZN(_00069_ ) );
BUF_X4 _23637_ ( .A(_08571_ ), .Z(_08573_ ) );
AOI21_X1 _23638_ ( .A(_08573_ ), .B1(_06080_ ), .B2(_06083_ ), .ZN(_00070_ ) );
NOR2_X1 _23639_ ( .A1(_06090_ ), .A2(_08572_ ), .ZN(_00071_ ) );
AOI21_X1 _23640_ ( .A(_08573_ ), .B1(_08568_ ), .B2(_06093_ ), .ZN(_00072_ ) );
NOR2_X1 _23641_ ( .A1(_06096_ ), .A2(_08572_ ), .ZN(_00073_ ) );
AOI21_X1 _23642_ ( .A(_08573_ ), .B1(_08568_ ), .B2(_06097_ ), .ZN(_00074_ ) );
NOR2_X1 _23643_ ( .A1(_06100_ ), .A2(_08572_ ), .ZN(_00075_ ) );
AOI21_X1 _23644_ ( .A(_08573_ ), .B1(_06104_ ), .B2(_06105_ ), .ZN(_00076_ ) );
NOR2_X1 _23645_ ( .A1(_06110_ ), .A2(_08572_ ), .ZN(_00077_ ) );
AOI21_X1 _23646_ ( .A(_08573_ ), .B1(_08568_ ), .B2(_06111_ ), .ZN(_00078_ ) );
AOI21_X1 _23647_ ( .A(_08573_ ), .B1(_08568_ ), .B2(_06112_ ), .ZN(_00079_ ) );
AOI21_X1 _23648_ ( .A(_08573_ ), .B1(_06114_ ), .B2(_06115_ ), .ZN(_00080_ ) );
NOR2_X1 _23649_ ( .A1(_06120_ ), .A2(_08572_ ), .ZN(_00081_ ) );
NOR2_X1 _23650_ ( .A1(_06123_ ), .A2(_08572_ ), .ZN(_00082_ ) );
NOR2_X1 _23651_ ( .A1(_06128_ ), .A2(_08572_ ), .ZN(_00083_ ) );
NOR2_X1 _23652_ ( .A1(_06132_ ), .A2(_08572_ ), .ZN(_00084_ ) );
BUF_X4 _23653_ ( .A(_08571_ ), .Z(_08574_ ) );
NOR2_X1 _23654_ ( .A1(_06136_ ), .A2(_08574_ ), .ZN(_00085_ ) );
NOR2_X1 _23655_ ( .A1(_06140_ ), .A2(_08574_ ), .ZN(_00086_ ) );
NOR2_X1 _23656_ ( .A1(_06669_ ), .A2(_08574_ ), .ZN(_00087_ ) );
NOR2_X1 _23657_ ( .A1(_07007_ ), .A2(_08574_ ), .ZN(_00088_ ) );
NOR2_X1 _23658_ ( .A1(_07315_ ), .A2(_08574_ ), .ZN(_00089_ ) );
NOR2_X1 _23659_ ( .A1(_07617_ ), .A2(_08574_ ), .ZN(_00090_ ) );
NOR2_X1 _23660_ ( .A1(_07913_ ), .A2(_08574_ ), .ZN(_00091_ ) );
AOI21_X1 _23661_ ( .A(_08573_ ), .B1(_07915_ ), .B2(_07916_ ), .ZN(_00092_ ) );
NOR2_X1 _23662_ ( .A1(_08228_ ), .A2(_08574_ ), .ZN(_00093_ ) );
AOI21_X1 _23663_ ( .A(_08573_ ), .B1(_08548_ ), .B2(_08549_ ), .ZN(_00094_ ) );
NOR2_X1 _23664_ ( .A1(_08554_ ), .A2(_08574_ ), .ZN(_00095_ ) );
AOI21_X1 _23665_ ( .A(_08573_ ), .B1(_06091_ ), .B2(_08555_ ), .ZN(_00096_ ) );
AOI21_X1 _23666_ ( .A(_08571_ ), .B1(_06091_ ), .B2(_08556_ ), .ZN(_00097_ ) );
AOI21_X1 _23667_ ( .A(_08571_ ), .B1(_06091_ ), .B2(_08557_ ), .ZN(_00098_ ) );
NOR2_X1 _23668_ ( .A1(_08562_ ), .A2(_08574_ ), .ZN(_00099_ ) );
AOI21_X1 _23669_ ( .A(_08571_ ), .B1(_06091_ ), .B2(_08563_ ), .ZN(_00100_ ) );
CLKBUF_X1 _23670_ ( .A(fanout_net_75 ), .Z(\u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _23671_ ( .A1(_08572_ ), .A2(_09110_ ), .ZN(\u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _23672_ ( .A1(_06075_ ), .A2(_09110_ ), .ZN(\u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _23673_ ( .A1(_08566_ ), .A2(_09110_ ), .ZN(\u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_E ) );
AND3_X1 _23674_ ( .A1(_08944_ ), .A2(_08920_ ), .A3(_08997_ ), .ZN(alu_result_out_$_XNOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__B_Y ) );
CLKGATE_X1 _23675_ ( .CK(clk ), .E(alu_result_out_$_XNOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__B_Y ), .GCK(_11608_ ) );
CLKGATE_X1 _23676_ ( .CK(clk ), .E(jump_en ), .GCK(_11609_ ) );
CLKGATE_X1 _23677_ ( .CK(clk ), .E(\u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_E ), .GCK(_11610_ ) );
CLKGATE_X1 _23678_ ( .CK(clk ), .E(\u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_E ), .GCK(_11611_ ) );
CLKGATE_X1 _23679_ ( .CK(clk ), .E(\u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_E ), .GCK(_11612_ ) );
CLKGATE_X1 _23680_ ( .CK(clk ), .E(\u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_E ), .GCK(_11613_ ) );
LOGIC0_X1 _23681_ ( .Z(_00000_ ) );
DFF_X1 ifu_rdata_$_SDFF_PP0__Q ( .D(_00001_ ), .CK(clk ), .Q(\ifu_rdata[2] ), .QN(alu_result_out_$_XNOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B_$_OR__Y_B_$_NOR__Y_A_$_XOR__Y_B_$_OR__Y_A_$_OR__Y_B ) );
DFF_X1 ifu_rdata_$_SDFF_PP0__Q_1 ( .D(_00002_ ), .CK(clk ), .Q(\ifu_rdata[0] ), .QN(_12019_ ) );
DFF_X1 ifu_rdata_$_SDFF_PP0__Q_2 ( .D(_00003_ ), .CK(clk ), .Q(\ifu_rdata[5] ), .QN(_12018_ ) );
DFF_X1 ifu_rdata_$_SDFF_PP0__Q_3 ( .D(_00004_ ), .CK(clk ), .Q(\ifu_rdata[4] ), .QN(_12017_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][31] ), .QN(_12020_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_1 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][30] ), .QN(_12016_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_10 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][21] ), .QN(_12015_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_11 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][20] ), .QN(_12014_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_12 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][19] ), .QN(_12013_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_13 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][18] ), .QN(_12012_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_14 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][17] ), .QN(_12011_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_15 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][16] ), .QN(_12010_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_16 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][15] ), .QN(_12009_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_17 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][14] ), .QN(_12008_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_18 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][13] ), .QN(_12007_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_19 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][12] ), .QN(_12006_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_2 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][29] ), .QN(_12005_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_20 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][11] ), .QN(_12004_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_21 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][10] ), .QN(_12003_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_22 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][9] ), .QN(_12002_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_23 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][8] ), .QN(_12001_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_24 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][7] ), .QN(_12000_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_25 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][6] ), .QN(_11999_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_26 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][5] ), .QN(_11998_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_27 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][4] ), .QN(_11997_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_28 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][3] ), .QN(_11996_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_29 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][2] ), .QN(_11995_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_3 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][28] ), .QN(_11994_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_30 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][1] ), .QN(_11993_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_31 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][0] ), .QN(_11992_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_4 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][27] ), .QN(_11991_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_5 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][26] ), .QN(_11990_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_6 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][25] ), .QN(_11989_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_7 ( .D(fanout_net_1 ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][24] ), .QN(_11988_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_8 ( .D(_00000_ ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][23] ), .QN(_11987_ ) );
DFF_X1 \u_gpr.regfile[0]_$_SDFFCE_PN0P__Q_9 ( .D(_00000_ ), .CK(_11613_ ), .Q(\u_gpr.regfile[0][22] ), .QN(_11986_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q ( .D(_00005_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][31] ), .QN(_11985_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_1 ( .D(_00006_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][30] ), .QN(_11984_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_10 ( .D(_00007_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][21] ), .QN(_11983_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_11 ( .D(_00008_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][20] ), .QN(_11982_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_12 ( .D(_00009_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][19] ), .QN(_11981_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_13 ( .D(_00010_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][18] ), .QN(_11980_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_14 ( .D(_00011_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][17] ), .QN(_11979_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_15 ( .D(_00012_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][16] ), .QN(_11978_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_16 ( .D(_00013_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][15] ), .QN(_11977_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_17 ( .D(_00014_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][14] ), .QN(_11976_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_18 ( .D(_00015_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][13] ), .QN(_11975_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_19 ( .D(_00016_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][12] ), .QN(_11974_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_2 ( .D(_00017_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][29] ), .QN(_11973_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_20 ( .D(_00018_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][11] ), .QN(_11972_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_21 ( .D(_00019_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][10] ), .QN(_11971_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_22 ( .D(_00020_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][9] ), .QN(_11970_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_23 ( .D(_00021_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][8] ), .QN(_11969_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_24 ( .D(_00022_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][7] ), .QN(_11968_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_25 ( .D(_00023_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][6] ), .QN(_11967_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_26 ( .D(_00024_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][5] ), .QN(_11966_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_27 ( .D(_00025_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][4] ), .QN(_11965_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_28 ( .D(_00026_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][3] ), .QN(_11964_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_29 ( .D(_00027_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][2] ), .QN(_11963_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_3 ( .D(_00028_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][28] ), .QN(_11962_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_30 ( .D(_00029_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][1] ), .QN(_11961_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_31 ( .D(_00030_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][0] ), .QN(_11960_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_4 ( .D(_00031_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][27] ), .QN(_11959_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_5 ( .D(_00032_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][26] ), .QN(_11958_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_6 ( .D(_00033_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][25] ), .QN(_11957_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_7 ( .D(_00034_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][24] ), .QN(_11956_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_8 ( .D(_00035_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][23] ), .QN(_11955_ ) );
DFF_X1 \u_gpr.regfile[1]_$_SDFFCE_PN0P__Q_9 ( .D(_00036_ ), .CK(_11612_ ), .Q(\u_gpr.regfile[1][22] ), .QN(_11954_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q ( .D(_00037_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][31] ), .QN(_11953_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_1 ( .D(_00038_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][30] ), .QN(_11952_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_10 ( .D(_00039_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][21] ), .QN(_11951_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_11 ( .D(_00040_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][20] ), .QN(_11950_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_12 ( .D(_00041_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][19] ), .QN(_11949_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_13 ( .D(_00042_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][18] ), .QN(_11948_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_14 ( .D(_00043_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][17] ), .QN(_11947_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_15 ( .D(_00044_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][16] ), .QN(_11946_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_16 ( .D(_00045_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][15] ), .QN(_11945_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_17 ( .D(_00046_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][14] ), .QN(_11944_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_18 ( .D(_00047_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][13] ), .QN(_11943_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_19 ( .D(_00048_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][12] ), .QN(_11942_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_2 ( .D(_00049_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][29] ), .QN(_11941_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_20 ( .D(_00050_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][11] ), .QN(_11940_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_21 ( .D(_00051_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][10] ), .QN(_11939_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_22 ( .D(_00052_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][9] ), .QN(_11938_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_23 ( .D(_00053_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][8] ), .QN(_11937_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_24 ( .D(_00054_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][7] ), .QN(_11936_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_25 ( .D(_00055_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][6] ), .QN(_11935_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_26 ( .D(_00056_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][5] ), .QN(_11934_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_27 ( .D(_00057_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][4] ), .QN(_11933_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_28 ( .D(_00058_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][3] ), .QN(_11932_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_29 ( .D(_00059_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][2] ), .QN(_11931_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_3 ( .D(_00060_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][28] ), .QN(_11930_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_30 ( .D(_00061_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][1] ), .QN(_11929_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_31 ( .D(_00062_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][0] ), .QN(_11928_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_4 ( .D(_00063_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][27] ), .QN(_11927_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_5 ( .D(_00064_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][26] ), .QN(_11926_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_6 ( .D(_00065_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][25] ), .QN(_11925_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_7 ( .D(_00066_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][24] ), .QN(_11924_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_8 ( .D(_00067_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][23] ), .QN(_11923_ ) );
DFF_X1 \u_gpr.regfile[2]_$_SDFFCE_PN0P__Q_9 ( .D(_00068_ ), .CK(_11611_ ), .Q(\u_gpr.regfile[2][22] ), .QN(_11922_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q ( .D(_00069_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][31] ), .QN(_11921_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_1 ( .D(_00070_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][30] ), .QN(_11920_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_10 ( .D(_00071_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][21] ), .QN(_11919_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_11 ( .D(_00072_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][20] ), .QN(_11918_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_12 ( .D(_00073_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][19] ), .QN(_11917_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_13 ( .D(_00074_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][18] ), .QN(_11916_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_14 ( .D(_00075_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][17] ), .QN(_11915_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_15 ( .D(_00076_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][16] ), .QN(_11914_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_16 ( .D(_00077_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][15] ), .QN(_11913_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_17 ( .D(_00078_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][14] ), .QN(_11912_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_18 ( .D(_00079_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][13] ), .QN(_11911_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_19 ( .D(_00080_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][12] ), .QN(_11910_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_2 ( .D(_00081_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][29] ), .QN(_11909_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_20 ( .D(_00082_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][11] ), .QN(_11908_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_21 ( .D(_00083_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][10] ), .QN(_11907_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_22 ( .D(_00084_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][9] ), .QN(_11906_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_23 ( .D(_00085_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][8] ), .QN(_11905_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_24 ( .D(_00086_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][7] ), .QN(_11904_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_25 ( .D(_00087_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][6] ), .QN(_11903_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_26 ( .D(_00088_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][5] ), .QN(_11902_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_27 ( .D(_00089_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][4] ), .QN(_11901_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_28 ( .D(_00090_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][3] ), .QN(_11900_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_29 ( .D(_00091_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][2] ), .QN(_11899_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_3 ( .D(_00092_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][28] ), .QN(_11898_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_30 ( .D(_00093_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][1] ), .QN(_11897_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_31 ( .D(_00094_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][0] ), .QN(_11896_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_4 ( .D(_00095_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][27] ), .QN(_11895_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_5 ( .D(_00096_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][26] ), .QN(_11894_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_6 ( .D(_00097_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][25] ), .QN(_11893_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_7 ( .D(_00098_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][24] ), .QN(_11892_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_8 ( .D(_00099_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][23] ), .QN(_11891_ ) );
DFF_X1 \u_gpr.regfile[3]_$_SDFFCE_PN0P__Q_9 ( .D(_00100_ ), .CK(_11610_ ), .Q(\u_gpr.regfile[3][22] ), .QN(_11890_ ) );
DFF_X1 \u_idu.inst_$_SDFF_PP0__Q ( .D(_00102_ ), .CK(clk ), .Q(\ifu_rdata[16] ), .QN(alu_result_out_$_XNOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B_$_OR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \u_idu.inst_$_SDFF_PP0__Q_1 ( .D(_00103_ ), .CK(clk ), .Q(\ifu_rdata[15] ), .QN(_11889_ ) );
DFF_X1 \u_idu.inst_$_SDFF_PP0__Q_2 ( .D(_00104_ ), .CK(clk ), .Q(\ifu_rdata[21] ), .QN(\u_ifu.jump_en_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_NOR__Y_A_$_OR__Y_B ) );
DFF_X1 \u_idu.inst_$_SDFF_PP0__Q_3 ( .D(_00105_ ), .CK(clk ), .Q(\ifu_rdata[20] ), .QN(alu_result_out_$_XNOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B_$_ORNOT__B_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \u_idu.inst_$_SDFF_PP0__Q_4 ( .D(_00106_ ), .CK(clk ), .Q(\ifu_rdata[8] ), .QN(_11888_ ) );
DFF_X1 \u_idu.inst_$_SDFF_PP0__Q_5 ( .D(_00107_ ), .CK(clk ), .Q(\ifu_rdata[7] ), .QN(_11887_ ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0P__Q ( .D(_00101_ ), .CK(_11609_ ), .Q(\pc_out[1] ), .QN(\u_gpr.gpr_wdata_$_ANDNOT__Y_30_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \u_ifu.pc_$_SDFFE_PP0P__Q_1 ( .D(_00108_ ), .CK(_11609_ ), .Q(\pc_out[0] ), .QN(_11886_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q ( .D(_00110_ ), .CK(clk ), .Q(\pc_out[30] ), .QN(dnpc_$_MUX__Y_1_A_$_NOT__Y_A_$_XOR__Y_B ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_1 ( .D(_00111_ ), .CK(clk ), .Q(\pc_out[29] ), .QN(_11885_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_10 ( .D(_00112_ ), .CK(clk ), .Q(\pc_out[20] ), .QN(dnpc_$_MUX__Y_11_A_$_NOT__Y_A_$_XOR__Y_B ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_11 ( .D(_00113_ ), .CK(clk ), .Q(\pc_out[19] ), .QN(_11884_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_12 ( .D(_00114_ ), .CK(clk ), .Q(\pc_out[18] ), .QN(dnpc_$_MUX__Y_13_A_$_NOT__Y_A_$_XOR__Y_B ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_13 ( .D(_00115_ ), .CK(clk ), .Q(\pc_out[17] ), .QN(_11883_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_14 ( .D(_00116_ ), .CK(clk ), .Q(\pc_out[16] ), .QN(dnpc_$_MUX__Y_15_A_$_NOT__Y_A_$_XOR__Y_B ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_15 ( .D(_00117_ ), .CK(clk ), .Q(\pc_out[15] ), .QN(_11882_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_16 ( .D(_00118_ ), .CK(clk ), .Q(\pc_out[14] ), .QN(dnpc_$_MUX__Y_17_A_$_NOT__Y_A_$_XOR__Y_B ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_17 ( .D(_00119_ ), .CK(clk ), .Q(\pc_out[13] ), .QN(_11881_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_18 ( .D(_00120_ ), .CK(clk ), .Q(\pc_out[12] ), .QN(_11880_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_19 ( .D(_00121_ ), .CK(clk ), .Q(\pc_out[11] ), .QN(_11879_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_2 ( .D(_00122_ ), .CK(clk ), .Q(\pc_out[28] ), .QN(dnpc_$_MUX__Y_3_A_$_NOT__Y_A_$_XOR__Y_B ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_20 ( .D(_00123_ ), .CK(clk ), .Q(\pc_out[10] ), .QN(dnpc_$_MUX__Y_21_A_$_NOT__Y_A_$_XOR__Y_B ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_21 ( .D(_00124_ ), .CK(clk ), .Q(\pc_out[9] ), .QN(_11878_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_22 ( .D(_00125_ ), .CK(clk ), .Q(\pc_out[8] ), .QN(dnpc_$_NOT__Y_1_A_$_MUX__Y_A_$_XOR__Y_B ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_23 ( .D(_00126_ ), .CK(clk ), .Q(\pc_out[7] ), .QN(_11877_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_24 ( .D(_00127_ ), .CK(clk ), .Q(\pc_out[6] ), .QN(dnpc_$_NOT__Y_3_A_$_MUX__Y_A_$_XOR__Y_B ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_25 ( .D(_00128_ ), .CK(clk ), .Q(\pc_out[5] ), .QN(_11876_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_26 ( .D(_00129_ ), .CK(clk ), .Q(\pc_out[4] ), .QN(dnpc_$_NOT__Y_5_A_$_MUX__Y_A_$_XOR__Y_B ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_27 ( .D(_00130_ ), .CK(clk ), .Q(\pc_out[3] ), .QN(_11875_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_28 ( .D(_00131_ ), .CK(clk ), .Q(\pc_out[2] ), .QN(dnpc_$_MUX__Y_22_A ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_3 ( .D(_00132_ ), .CK(clk ), .Q(\pc_out[27] ), .QN(_11874_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_4 ( .D(_00133_ ), .CK(clk ), .Q(\pc_out[26] ), .QN(dnpc_$_MUX__Y_5_A_$_NOT__Y_A_$_XOR__Y_B ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_5 ( .D(_00134_ ), .CK(clk ), .Q(\pc_out[25] ), .QN(_11873_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_6 ( .D(_00135_ ), .CK(clk ), .Q(\pc_out[24] ), .QN(_11872_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_7 ( .D(_00136_ ), .CK(clk ), .Q(\pc_out[23] ), .QN(_11871_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_8 ( .D(_00137_ ), .CK(clk ), .Q(\pc_out[22] ), .QN(dnpc_$_MUX__Y_9_A_$_NOT__Y_A_$_XOR__Y_B ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_9 ( .D(_00138_ ), .CK(clk ), .Q(\pc_out[21] ), .QN(_11870_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP1__Q ( .D(_00139_ ), .CK(clk ), .Q(\pc_out[31] ), .QN(_12021_ ) );
DFF_X1 \u_ifu.reset_sync_$_DFF_P__Q ( .D(fanout_net_75 ), .CK(clk ), .Q(\u_ifu.reset_sync ), .QN(dnpc_$_NOT__Y_A_$_ANDNOT__B_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q ( .D(_00109_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4388] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1 ( .D(_00140_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4387] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_10 ( .D(_00141_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4354] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_100 ( .D(_00142_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4000] ), .QN(_11869_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1000 ( .D(_00143_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[388] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1001 ( .D(_00144_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[387] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1002 ( .D(_00145_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[386] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1003 ( .D(_00146_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[385] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1004 ( .D(_00147_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[384] ), .QN(_11868_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1005 ( .D(_00148_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[359] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1006 ( .D(_00149_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[358] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1007 ( .D(_00150_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[357] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1008 ( .D(_00151_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[356] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1009 ( .D(_00152_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[355] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_101 ( .D(_00153_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3975] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1010 ( .D(_00154_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[354] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1011 ( .D(_00155_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[353] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1012 ( .D(_00156_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[352] ), .QN(_11867_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1013 ( .D(_00157_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[327] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1014 ( .D(_00158_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[326] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1015 ( .D(_00159_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[325] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1016 ( .D(_00160_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[324] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1017 ( .D(_00161_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[323] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1018 ( .D(_00162_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[322] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1019 ( .D(_00163_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[321] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_102 ( .D(_00164_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3974] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1020 ( .D(_00165_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[320] ), .QN(_11866_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1021 ( .D(_00166_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[295] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1022 ( .D(_00167_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[294] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1023 ( .D(_00168_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[293] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1024 ( .D(_00169_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[292] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1025 ( .D(_00170_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[291] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1026 ( .D(_00171_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[290] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1027 ( .D(_00172_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[289] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1028 ( .D(_00173_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[288] ), .QN(_11865_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1029 ( .D(_00174_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[263] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_103 ( .D(_00175_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3973] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1030 ( .D(_00176_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[262] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1031 ( .D(_00177_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[261] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1032 ( .D(_00178_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[260] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1033 ( .D(_00179_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[259] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1034 ( .D(_00180_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[258] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1035 ( .D(_00181_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[257] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1036 ( .D(_00182_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[256] ), .QN(_11864_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1037 ( .D(_00183_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[231] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1038 ( .D(_00184_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[230] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1039 ( .D(_00185_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[229] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_104 ( .D(_00186_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3972] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1040 ( .D(_00187_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[228] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1041 ( .D(_00188_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[227] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1042 ( .D(_00189_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[226] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1043 ( .D(_00190_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[225] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1044 ( .D(_00191_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[224] ), .QN(_11863_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1045 ( .D(_00192_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[199] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1046 ( .D(_00193_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[198] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1047 ( .D(_00194_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[197] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1048 ( .D(_00195_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[196] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1049 ( .D(_00196_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[195] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_105 ( .D(_00197_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3971] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1050 ( .D(_00198_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[194] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1051 ( .D(_00199_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[193] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1052 ( .D(_00200_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[192] ), .QN(_11862_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1053 ( .D(_00201_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[167] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1054 ( .D(_00202_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[166] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1055 ( .D(_00203_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[165] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1056 ( .D(_00204_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[164] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1057 ( .D(_00205_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[163] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1058 ( .D(_00206_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[162] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1059 ( .D(_00207_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[161] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_106 ( .D(_00208_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3970] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1060 ( .D(_00209_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[160] ), .QN(_11861_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1061 ( .D(_00210_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[135] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1062 ( .D(_00211_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[134] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1063 ( .D(_00212_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[133] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1064 ( .D(_00213_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[132] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1065 ( .D(_00214_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[131] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1066 ( .D(_00215_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[130] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1067 ( .D(_00216_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[129] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1068 ( .D(_00217_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[128] ), .QN(_11860_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1069 ( .D(_00218_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[103] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_107 ( .D(_00219_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3969] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1070 ( .D(_00220_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[102] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1071 ( .D(_00221_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[101] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1072 ( .D(_00222_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[100] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1073 ( .D(_00223_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[99] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1074 ( .D(_00224_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[98] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1075 ( .D(_00225_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[97] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1076 ( .D(_00226_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[96] ), .QN(_11859_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1077 ( .D(_00227_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[71] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1078 ( .D(_00228_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[70] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1079 ( .D(_00229_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[69] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_108 ( .D(_00230_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3968] ), .QN(_11858_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1080 ( .D(_00231_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[68] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1081 ( .D(_00232_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[67] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1082 ( .D(_00233_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[66] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1083 ( .D(_00234_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[65] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1084 ( .D(_00235_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[64] ), .QN(_11857_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1085 ( .D(_00236_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[39] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1086 ( .D(_00237_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[38] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1087 ( .D(_00238_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[37] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1088 ( .D(_00239_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[36] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1089 ( .D(_00240_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[35] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_109 ( .D(_00241_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3943] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1090 ( .D(_00242_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[34] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1091 ( .D(_00243_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[33] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1092 ( .D(_00244_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[32] ), .QN(_11856_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1093 ( .D(_00245_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1094 ( .D(_00246_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1095 ( .D(_00247_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1096 ( .D(_00248_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1097 ( .D(_00249_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1098 ( .D(_00250_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1099 ( .D(_00251_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_11 ( .D(_00252_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4353] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_110 ( .D(_00253_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3942] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1100 ( .D(_00254_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[0] ), .QN(_11855_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1101 ( .D(_00255_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8167] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1102 ( .D(_00256_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8166] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1103 ( .D(_00257_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8165] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1104 ( .D(_00258_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8164] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1105 ( .D(_00259_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8163] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1106 ( .D(_00260_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8162] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1107 ( .D(_00261_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8161] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1108 ( .D(_00262_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8160] ), .QN(_11854_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1109 ( .D(_00263_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8135] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_111 ( .D(_00264_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3941] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1110 ( .D(_00265_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8134] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1111 ( .D(_00266_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8133] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1112 ( .D(_00267_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8132] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1113 ( .D(_00268_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8131] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1114 ( .D(_00269_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8130] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1115 ( .D(_00270_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8129] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1116 ( .D(_00271_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8128] ), .QN(_11853_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1117 ( .D(_00272_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8103] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1118 ( .D(_00273_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8102] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1119 ( .D(_00274_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8101] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_112 ( .D(_00275_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3940] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1120 ( .D(_00276_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8100] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1121 ( .D(_00277_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8099] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1122 ( .D(_00278_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8098] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1123 ( .D(_00279_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8097] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1124 ( .D(_00280_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8096] ), .QN(_11852_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1125 ( .D(_00281_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8071] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1126 ( .D(_00282_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8070] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1127 ( .D(_00283_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8069] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1128 ( .D(_00284_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8068] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1129 ( .D(_00285_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8067] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_113 ( .D(_00286_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3939] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1130 ( .D(_00287_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8066] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1131 ( .D(_00288_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8065] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1132 ( .D(_00289_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8064] ), .QN(_11851_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1133 ( .D(_00290_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8039] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1134 ( .D(_00291_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8038] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1135 ( .D(_00292_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8037] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1136 ( .D(_00293_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8036] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1137 ( .D(_00294_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8035] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1138 ( .D(_00295_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8034] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1139 ( .D(_00296_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8033] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_114 ( .D(_00297_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3938] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1140 ( .D(_00298_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8032] ), .QN(_11850_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1141 ( .D(_00299_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8007] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1142 ( .D(_00300_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8006] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1143 ( .D(_00301_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8005] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1144 ( .D(_00302_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8004] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1145 ( .D(_00303_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8003] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1146 ( .D(_00304_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8002] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1147 ( .D(_00305_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8001] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1148 ( .D(_00306_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[8000] ), .QN(_11849_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1149 ( .D(_00307_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7975] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_115 ( .D(_00308_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3937] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1150 ( .D(_00309_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7974] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1151 ( .D(_00310_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7973] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1152 ( .D(_00311_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7972] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1153 ( .D(_00312_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7971] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1154 ( .D(_00313_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7970] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1155 ( .D(_00314_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7969] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1156 ( .D(_00315_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7968] ), .QN(_11848_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1157 ( .D(_00316_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7943] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1158 ( .D(_00317_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7942] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1159 ( .D(_00318_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7941] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_116 ( .D(_00319_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3936] ), .QN(_11847_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1160 ( .D(_00320_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7940] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1161 ( .D(_00321_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7939] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1162 ( .D(_00322_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7938] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1163 ( .D(_00323_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7937] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1164 ( .D(_00324_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7936] ), .QN(_11846_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1165 ( .D(_00325_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7911] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1166 ( .D(_00326_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7910] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1167 ( .D(_00327_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7909] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1168 ( .D(_00328_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7908] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1169 ( .D(_00329_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7907] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_117 ( .D(_00330_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3911] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1170 ( .D(_00331_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7906] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1171 ( .D(_00332_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7905] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1172 ( .D(_00333_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7904] ), .QN(_11845_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1173 ( .D(_00334_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7879] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1174 ( .D(_00335_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7878] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1175 ( .D(_00336_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7877] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1176 ( .D(_00337_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7876] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1177 ( .D(_00338_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7875] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1178 ( .D(_00339_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7874] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1179 ( .D(_00340_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7873] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_118 ( .D(_00341_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3910] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1180 ( .D(_00342_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7872] ), .QN(_11844_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1181 ( .D(_00343_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7847] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1182 ( .D(_00344_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7846] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1183 ( .D(_00345_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7845] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1184 ( .D(_00346_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7844] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1185 ( .D(_00347_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7843] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1186 ( .D(_00348_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7842] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1187 ( .D(_00349_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7841] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1188 ( .D(_00350_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7840] ), .QN(_11843_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1189 ( .D(_00351_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7815] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_119 ( .D(_00352_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3909] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1190 ( .D(_00353_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7814] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1191 ( .D(_00354_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7813] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1192 ( .D(_00355_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7812] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1193 ( .D(_00356_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7811] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1194 ( .D(_00357_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7810] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1195 ( .D(_00358_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7809] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1196 ( .D(_00359_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7808] ), .QN(_11842_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1197 ( .D(_00360_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7783] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1198 ( .D(_00361_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7782] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1199 ( .D(_00362_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7781] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_12 ( .D(_00363_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4352] ), .QN(_11841_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_120 ( .D(_00364_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3908] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1200 ( .D(_00365_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7780] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1201 ( .D(_00366_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7779] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1202 ( .D(_00367_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7778] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1203 ( .D(_00368_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7777] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1204 ( .D(_00369_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7776] ), .QN(_11840_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1205 ( .D(_00370_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7751] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1206 ( .D(_00371_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7750] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1207 ( .D(_00372_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7749] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1208 ( .D(_00373_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7748] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1209 ( .D(_00374_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7747] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_121 ( .D(_00375_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3907] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1210 ( .D(_00376_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7746] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1211 ( .D(_00377_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7745] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1212 ( .D(_00378_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7744] ), .QN(_11839_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1213 ( .D(_00379_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7719] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1214 ( .D(_00380_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7718] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1215 ( .D(_00381_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7717] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1216 ( .D(_00382_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7716] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1217 ( .D(_00383_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7715] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1218 ( .D(_00384_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7714] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1219 ( .D(_00385_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7713] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_122 ( .D(_00386_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3906] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1220 ( .D(_00387_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7712] ), .QN(_11838_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1221 ( .D(_00388_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7687] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1222 ( .D(_00389_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7686] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1223 ( .D(_00390_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7685] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1224 ( .D(_00391_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7684] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1225 ( .D(_00392_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7683] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1226 ( .D(_00393_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7682] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1227 ( .D(_00394_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7681] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1228 ( .D(_00395_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7680] ), .QN(_11837_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1229 ( .D(_00396_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7655] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_123 ( .D(_00397_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3905] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1230 ( .D(_00398_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7654] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1231 ( .D(_00399_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7653] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1232 ( .D(_00400_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7652] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1233 ( .D(_00401_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7651] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1234 ( .D(_00402_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7650] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1235 ( .D(_00403_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7649] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1236 ( .D(_00404_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7648] ), .QN(_11836_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1237 ( .D(_00405_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7623] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1238 ( .D(_00406_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7622] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1239 ( .D(_00407_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7621] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_124 ( .D(_00408_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3904] ), .QN(_11835_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1240 ( .D(_00409_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7620] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1241 ( .D(_00410_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7619] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1242 ( .D(_00411_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7618] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1243 ( .D(_00412_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7617] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1244 ( .D(_00413_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7616] ), .QN(_11834_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1245 ( .D(_00414_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7591] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1246 ( .D(_00415_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7590] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1247 ( .D(_00416_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7589] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1248 ( .D(_00417_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7588] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1249 ( .D(_00418_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7587] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_125 ( .D(_00419_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3879] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1250 ( .D(_00420_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7586] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1251 ( .D(_00421_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7585] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1252 ( .D(_00422_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7584] ), .QN(_11833_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1253 ( .D(_00423_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7559] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1254 ( .D(_00424_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7558] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1255 ( .D(_00425_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7557] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1256 ( .D(_00426_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7556] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1257 ( .D(_00427_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7555] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1258 ( .D(_00428_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7554] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1259 ( .D(_00429_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7553] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_126 ( .D(_00430_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3878] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1260 ( .D(_00431_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7552] ), .QN(_11832_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1261 ( .D(_00432_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7527] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1262 ( .D(_00433_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7526] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1263 ( .D(_00434_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7525] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1264 ( .D(_00435_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7524] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1265 ( .D(_00436_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7523] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1266 ( .D(_00437_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7522] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1267 ( .D(_00438_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7521] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1268 ( .D(_00439_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7520] ), .QN(_11831_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1269 ( .D(_00440_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7495] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_127 ( .D(_00441_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3877] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1270 ( .D(_00442_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7494] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1271 ( .D(_00443_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7493] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1272 ( .D(_00444_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7492] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1273 ( .D(_00445_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7491] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1274 ( .D(_00446_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7490] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1275 ( .D(_00447_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7489] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1276 ( .D(_00448_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7488] ), .QN(_11830_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1277 ( .D(_00449_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7463] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1278 ( .D(_00450_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7462] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1279 ( .D(_00451_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7461] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_128 ( .D(_00452_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3876] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1280 ( .D(_00453_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7460] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1281 ( .D(_00454_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7459] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1282 ( .D(_00455_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7458] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1283 ( .D(_00456_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7457] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1284 ( .D(_00457_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7456] ), .QN(_11829_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1285 ( .D(_00458_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7431] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1286 ( .D(_00459_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7430] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1287 ( .D(_00460_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7429] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1288 ( .D(_00461_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7428] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1289 ( .D(_00462_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7427] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_129 ( .D(_00463_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3875] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1290 ( .D(_00464_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7426] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1291 ( .D(_00465_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7425] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1292 ( .D(_00466_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7424] ), .QN(_11828_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1293 ( .D(_00467_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7399] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1294 ( .D(_00468_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7398] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1295 ( .D(_00469_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7397] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1296 ( .D(_00470_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7396] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1297 ( .D(_00471_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7395] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1298 ( .D(_00472_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7394] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1299 ( .D(_00473_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7393] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_13 ( .D(_00474_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4327] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_130 ( .D(_00475_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3874] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1300 ( .D(_00476_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7392] ), .QN(_11827_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1301 ( .D(_00477_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7367] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1302 ( .D(_00478_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7366] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1303 ( .D(_00479_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7365] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1304 ( .D(_00480_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7364] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1305 ( .D(_00481_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7363] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1306 ( .D(_00482_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7362] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1307 ( .D(_00483_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7361] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1308 ( .D(_00484_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7360] ), .QN(_11826_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1309 ( .D(_00485_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7335] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_131 ( .D(_00486_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3873] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1310 ( .D(_00487_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7334] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1311 ( .D(_00488_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7333] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1312 ( .D(_00489_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7332] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1313 ( .D(_00490_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7331] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1314 ( .D(_00491_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7330] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1315 ( .D(_00492_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7329] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1316 ( .D(_00493_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7328] ), .QN(_11825_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1317 ( .D(_00494_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7303] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1318 ( .D(_00495_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7302] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1319 ( .D(_00496_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7301] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_132 ( .D(_00497_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3872] ), .QN(_11824_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1320 ( .D(_00498_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7300] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1321 ( .D(_00499_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7299] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1322 ( .D(_00500_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7298] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1323 ( .D(_00501_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7297] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1324 ( .D(_00502_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7296] ), .QN(_11823_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1325 ( .D(_00503_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7271] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1326 ( .D(_00504_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7270] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1327 ( .D(_00505_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7269] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1328 ( .D(_00506_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7268] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1329 ( .D(_00507_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7267] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_133 ( .D(_00508_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3847] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1330 ( .D(_00509_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7266] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1331 ( .D(_00510_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7265] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1332 ( .D(_00511_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7264] ), .QN(_11822_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1333 ( .D(_00512_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7239] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1334 ( .D(_00513_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7238] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1335 ( .D(_00514_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7237] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1336 ( .D(_00515_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7236] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1337 ( .D(_00516_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7235] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1338 ( .D(_00517_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7234] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1339 ( .D(_00518_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7233] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_134 ( .D(_00519_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3846] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1340 ( .D(_00520_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7232] ), .QN(_11821_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1341 ( .D(_00521_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7207] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1342 ( .D(_00522_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7206] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1343 ( .D(_00523_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7205] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1344 ( .D(_00524_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7204] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1345 ( .D(_00525_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7203] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1346 ( .D(_00526_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7202] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1347 ( .D(_00527_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7201] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1348 ( .D(_00528_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7200] ), .QN(_11820_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1349 ( .D(_00529_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7175] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_135 ( .D(_00530_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3845] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1350 ( .D(_00531_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7174] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1351 ( .D(_00532_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7173] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1352 ( .D(_00533_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7172] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1353 ( .D(_00534_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7171] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1354 ( .D(_00535_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7170] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1355 ( .D(_00536_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7169] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1356 ( .D(_00537_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7168] ), .QN(_11819_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1357 ( .D(_00538_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7143] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1358 ( .D(_00539_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7142] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1359 ( .D(_00540_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7141] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_136 ( .D(_00541_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3844] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1360 ( .D(_00542_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7140] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1361 ( .D(_00543_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7139] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1362 ( .D(_00544_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7138] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1363 ( .D(_00545_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7137] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1364 ( .D(_00546_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7136] ), .QN(_11818_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1365 ( .D(_00547_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7111] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1366 ( .D(_00548_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7110] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1367 ( .D(_00549_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7109] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1368 ( .D(_00550_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7108] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1369 ( .D(_00551_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7107] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_137 ( .D(_00552_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3843] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1370 ( .D(_00553_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7106] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1371 ( .D(_00554_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7105] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1372 ( .D(_00555_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7104] ), .QN(_11817_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1373 ( .D(_00556_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7079] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1374 ( .D(_00557_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7078] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1375 ( .D(_00558_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7077] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1376 ( .D(_00559_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7076] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1377 ( .D(_00560_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7075] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1378 ( .D(_00561_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7074] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1379 ( .D(_00562_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7073] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_138 ( .D(_00563_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3842] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1380 ( .D(_00564_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7072] ), .QN(_11816_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1381 ( .D(_00565_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7047] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1382 ( .D(_00566_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7046] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1383 ( .D(_00567_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7045] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1384 ( .D(_00568_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7044] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1385 ( .D(_00569_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7043] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1386 ( .D(_00570_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7042] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1387 ( .D(_00571_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7041] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1388 ( .D(_00572_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7040] ), .QN(_11815_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1389 ( .D(_00573_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7015] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_139 ( .D(_00574_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3841] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1390 ( .D(_00575_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7014] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1391 ( .D(_00576_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7013] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1392 ( .D(_00577_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7012] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1393 ( .D(_00578_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7011] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1394 ( .D(_00579_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7010] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1395 ( .D(_00580_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7009] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1396 ( .D(_00581_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[7008] ), .QN(_11814_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1397 ( .D(_00582_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6983] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1398 ( .D(_00583_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6982] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1399 ( .D(_00584_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6981] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_14 ( .D(_00585_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4326] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_140 ( .D(_00586_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3840] ), .QN(_11813_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1400 ( .D(_00587_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6980] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1401 ( .D(_00588_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6979] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1402 ( .D(_00589_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6978] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1403 ( .D(_00590_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6977] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1404 ( .D(_00591_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6976] ), .QN(_11812_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1405 ( .D(_00592_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6951] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1406 ( .D(_00593_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6950] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1407 ( .D(_00594_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6949] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1408 ( .D(_00595_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6948] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1409 ( .D(_00596_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6947] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_141 ( .D(_00597_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3815] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1410 ( .D(_00598_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6946] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1411 ( .D(_00599_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6945] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1412 ( .D(_00600_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6944] ), .QN(_11811_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1413 ( .D(_00601_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6919] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1414 ( .D(_00602_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6918] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1415 ( .D(_00603_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6917] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1416 ( .D(_00604_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6916] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1417 ( .D(_00605_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6915] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1418 ( .D(_00606_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6914] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1419 ( .D(_00607_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6913] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_142 ( .D(_00608_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3814] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1420 ( .D(_00609_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6912] ), .QN(_11810_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1421 ( .D(_00610_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6887] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1422 ( .D(_00611_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6886] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1423 ( .D(_00612_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6885] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1424 ( .D(_00613_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6884] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1425 ( .D(_00614_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6883] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1426 ( .D(_00615_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6882] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1427 ( .D(_00616_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6881] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1428 ( .D(_00617_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6880] ), .QN(_11809_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1429 ( .D(_00618_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6855] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_143 ( .D(_00619_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3813] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1430 ( .D(_00620_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6854] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1431 ( .D(_00621_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6853] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1432 ( .D(_00622_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6852] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1433 ( .D(_00623_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6851] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1434 ( .D(_00624_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6850] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1435 ( .D(_00625_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6849] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1436 ( .D(_00626_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6848] ), .QN(_11808_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1437 ( .D(_00627_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6823] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1438 ( .D(_00628_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6822] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1439 ( .D(_00629_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6821] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_144 ( .D(_00630_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3812] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1440 ( .D(_00631_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6820] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1441 ( .D(_00632_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6819] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1442 ( .D(_00633_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6818] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1443 ( .D(_00634_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6817] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1444 ( .D(_00635_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6816] ), .QN(_11807_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1445 ( .D(_00636_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6791] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1446 ( .D(_00637_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6790] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1447 ( .D(_00638_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6789] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1448 ( .D(_00639_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6788] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1449 ( .D(_00640_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6787] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_145 ( .D(_00641_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3811] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1450 ( .D(_00642_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6786] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1451 ( .D(_00643_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6785] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1452 ( .D(_00644_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6784] ), .QN(_11806_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1453 ( .D(_00645_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6759] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1454 ( .D(_00646_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6758] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1455 ( .D(_00647_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6757] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1456 ( .D(_00648_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6756] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1457 ( .D(_00649_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6755] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1458 ( .D(_00650_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6754] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1459 ( .D(_00651_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6753] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_146 ( .D(_00652_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3810] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1460 ( .D(_00653_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6752] ), .QN(_11805_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1461 ( .D(_00654_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6727] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1462 ( .D(_00655_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6726] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1463 ( .D(_00656_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6725] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1464 ( .D(_00657_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6724] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1465 ( .D(_00658_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6723] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1466 ( .D(_00659_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6722] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1467 ( .D(_00660_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6721] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1468 ( .D(_00661_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6720] ), .QN(_11804_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1469 ( .D(_00662_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6695] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_147 ( .D(_00663_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3809] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1470 ( .D(_00664_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6694] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1471 ( .D(_00665_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6693] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1472 ( .D(_00666_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6692] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1473 ( .D(_00667_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6691] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1474 ( .D(_00668_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6690] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1475 ( .D(_00669_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6689] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1476 ( .D(_00670_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6688] ), .QN(_11803_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1477 ( .D(_00671_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6663] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1478 ( .D(_00672_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6662] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1479 ( .D(_00673_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6661] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_148 ( .D(_00674_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3808] ), .QN(_11802_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1480 ( .D(_00675_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6660] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1481 ( .D(_00676_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6659] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1482 ( .D(_00677_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6658] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1483 ( .D(_00678_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6657] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1484 ( .D(_00679_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6656] ), .QN(_11801_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1485 ( .D(_00680_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6631] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1486 ( .D(_00681_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6630] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1487 ( .D(_00682_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6629] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1488 ( .D(_00683_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6628] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1489 ( .D(_00684_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6627] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_149 ( .D(_00685_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3783] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1490 ( .D(_00686_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6626] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1491 ( .D(_00687_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6625] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1492 ( .D(_00688_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6624] ), .QN(_11800_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1493 ( .D(_00689_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6599] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1494 ( .D(_00690_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6598] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1495 ( .D(_00691_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6597] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1496 ( .D(_00692_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6596] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1497 ( .D(_00693_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6595] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1498 ( .D(_00694_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6594] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1499 ( .D(_00695_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6593] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_15 ( .D(_00696_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4325] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_150 ( .D(_00697_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3782] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1500 ( .D(_00698_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6592] ), .QN(_11799_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1501 ( .D(_00699_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6567] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1502 ( .D(_00700_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6566] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1503 ( .D(_00701_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6565] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1504 ( .D(_00702_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6564] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1505 ( .D(_00703_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6563] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1506 ( .D(_00704_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6562] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1507 ( .D(_00705_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6561] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1508 ( .D(_00706_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6560] ), .QN(_11798_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1509 ( .D(_00707_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6535] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_151 ( .D(_00708_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3781] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1510 ( .D(_00709_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6534] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1511 ( .D(_00710_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6533] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1512 ( .D(_00711_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6532] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1513 ( .D(_00712_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6531] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1514 ( .D(_00713_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6530] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1515 ( .D(_00714_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6529] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1516 ( .D(_00715_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6528] ), .QN(_11797_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1517 ( .D(_00716_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6503] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1518 ( .D(_00717_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6502] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1519 ( .D(_00718_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6501] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_152 ( .D(_00719_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3780] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1520 ( .D(_00720_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6500] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1521 ( .D(_00721_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6499] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1522 ( .D(_00722_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6498] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1523 ( .D(_00723_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6497] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1524 ( .D(_00724_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6496] ), .QN(_11796_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1525 ( .D(_00725_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6471] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1526 ( .D(_00726_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6470] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1527 ( .D(_00727_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6469] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1528 ( .D(_00728_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6468] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1529 ( .D(_00729_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6467] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_153 ( .D(_00730_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3779] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1530 ( .D(_00731_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6466] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1531 ( .D(_00732_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6465] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1532 ( .D(_00733_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6464] ), .QN(_11795_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1533 ( .D(_00734_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6439] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1534 ( .D(_00735_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6438] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1535 ( .D(_00736_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6437] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1536 ( .D(_00737_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6436] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1537 ( .D(_00738_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6435] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1538 ( .D(_00739_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6434] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1539 ( .D(_00740_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6433] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_154 ( .D(_00741_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3778] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1540 ( .D(_00742_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6432] ), .QN(_11794_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1541 ( .D(_00743_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6407] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1542 ( .D(_00744_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6406] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1543 ( .D(_00745_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6405] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1544 ( .D(_00746_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6404] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1545 ( .D(_00747_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6403] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1546 ( .D(_00748_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6402] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1547 ( .D(_00749_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6401] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1548 ( .D(_00750_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6400] ), .QN(_11793_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1549 ( .D(_00751_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6375] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_155 ( .D(_00752_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3777] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1550 ( .D(_00753_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6374] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1551 ( .D(_00754_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6373] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1552 ( .D(_00755_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6372] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1553 ( .D(_00756_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6371] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1554 ( .D(_00757_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6370] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1555 ( .D(_00758_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6369] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1556 ( .D(_00759_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6368] ), .QN(_11792_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1557 ( .D(_00760_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6343] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1558 ( .D(_00761_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6342] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1559 ( .D(_00762_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6341] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_156 ( .D(_00763_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3776] ), .QN(_11791_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1560 ( .D(_00764_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6340] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1561 ( .D(_00765_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6339] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1562 ( .D(_00766_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6338] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1563 ( .D(_00767_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6337] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1564 ( .D(_00768_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6336] ), .QN(_11790_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1565 ( .D(_00769_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6311] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1566 ( .D(_00770_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6310] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1567 ( .D(_00771_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6309] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1568 ( .D(_00772_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6308] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1569 ( .D(_00773_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6307] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_157 ( .D(_00774_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3751] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1570 ( .D(_00775_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6306] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1571 ( .D(_00776_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6305] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1572 ( .D(_00777_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6304] ), .QN(_11789_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1573 ( .D(_00778_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6279] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1574 ( .D(_00779_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6278] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1575 ( .D(_00780_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6277] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1576 ( .D(_00781_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6276] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1577 ( .D(_00782_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6275] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1578 ( .D(_00783_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6274] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1579 ( .D(_00784_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6273] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_158 ( .D(_00785_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3750] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1580 ( .D(_00786_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6272] ), .QN(_11788_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1581 ( .D(_00787_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6247] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1582 ( .D(_00788_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6246] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1583 ( .D(_00789_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6245] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1584 ( .D(_00790_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6244] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1585 ( .D(_00791_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6243] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1586 ( .D(_00792_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6242] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1587 ( .D(_00793_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6241] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1588 ( .D(_00794_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6240] ), .QN(_11787_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1589 ( .D(_00795_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6215] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_159 ( .D(_00796_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3749] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1590 ( .D(_00797_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6214] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1591 ( .D(_00798_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6213] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1592 ( .D(_00799_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6212] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1593 ( .D(_00800_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6211] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1594 ( .D(_00801_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6210] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1595 ( .D(_00802_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6209] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1596 ( .D(_00803_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6208] ), .QN(_11786_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1597 ( .D(_00804_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6183] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1598 ( .D(_00805_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6182] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1599 ( .D(_00806_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6181] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_16 ( .D(_00807_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4324] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_160 ( .D(_00808_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3748] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1600 ( .D(_00809_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6180] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1601 ( .D(_00810_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6179] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1602 ( .D(_00811_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6178] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1603 ( .D(_00812_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6177] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1604 ( .D(_00813_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6176] ), .QN(_11785_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1605 ( .D(_00814_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6151] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1606 ( .D(_00815_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6150] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1607 ( .D(_00816_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6149] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1608 ( .D(_00817_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6148] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1609 ( .D(_00818_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6147] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_161 ( .D(_00819_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3747] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1610 ( .D(_00820_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6146] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1611 ( .D(_00821_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6145] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1612 ( .D(_00822_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6144] ), .QN(_11784_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1613 ( .D(_00823_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6119] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1614 ( .D(_00824_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6118] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1615 ( .D(_00825_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6117] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1616 ( .D(_00826_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6116] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1617 ( .D(_00827_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6115] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1618 ( .D(_00828_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6114] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1619 ( .D(_00829_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6113] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_162 ( .D(_00830_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3746] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1620 ( .D(_00831_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6112] ), .QN(_11783_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1621 ( .D(_00832_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6087] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1622 ( .D(_00833_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6086] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1623 ( .D(_00834_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6085] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1624 ( .D(_00835_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6084] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1625 ( .D(_00836_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6083] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1626 ( .D(_00837_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6082] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1627 ( .D(_00838_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6081] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1628 ( .D(_00839_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6080] ), .QN(_11782_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1629 ( .D(_00840_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6055] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_163 ( .D(_00841_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3745] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1630 ( .D(_00842_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6054] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1631 ( .D(_00843_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6053] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1632 ( .D(_00844_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6052] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1633 ( .D(_00845_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6051] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1634 ( .D(_00846_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6050] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1635 ( .D(_00847_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6049] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1636 ( .D(_00848_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6048] ), .QN(_11781_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1637 ( .D(_00849_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6023] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1638 ( .D(_00850_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6022] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1639 ( .D(_00851_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6021] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_164 ( .D(_00852_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3744] ), .QN(_11780_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1640 ( .D(_00853_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6020] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1641 ( .D(_00854_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6019] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1642 ( .D(_00855_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6018] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1643 ( .D(_00856_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6017] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1644 ( .D(_00857_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[6016] ), .QN(_11779_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1645 ( .D(_00858_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5991] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1646 ( .D(_00859_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5990] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1647 ( .D(_00860_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5989] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1648 ( .D(_00861_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5988] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1649 ( .D(_00862_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5987] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_165 ( .D(_00863_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3719] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1650 ( .D(_00864_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5986] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1651 ( .D(_00865_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5985] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1652 ( .D(_00866_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5984] ), .QN(_11778_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1653 ( .D(_00867_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5959] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1654 ( .D(_00868_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5958] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1655 ( .D(_00869_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5957] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1656 ( .D(_00870_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5956] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1657 ( .D(_00871_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5955] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1658 ( .D(_00872_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5954] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1659 ( .D(_00873_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5953] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_166 ( .D(_00874_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3718] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1660 ( .D(_00875_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5952] ), .QN(_11777_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1661 ( .D(_00876_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5927] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1662 ( .D(_00877_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5926] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1663 ( .D(_00878_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5925] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1664 ( .D(_00879_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5924] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1665 ( .D(_00880_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5923] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1666 ( .D(_00881_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5922] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1667 ( .D(_00882_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5921] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1668 ( .D(_00883_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5920] ), .QN(_11776_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1669 ( .D(_00884_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5895] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_167 ( .D(_00885_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3717] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1670 ( .D(_00886_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5894] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1671 ( .D(_00887_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5893] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1672 ( .D(_00888_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5892] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1673 ( .D(_00889_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5891] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1674 ( .D(_00890_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5890] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1675 ( .D(_00891_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5889] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1676 ( .D(_00892_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5888] ), .QN(_11775_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1677 ( .D(_00893_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5863] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1678 ( .D(_00894_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5862] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1679 ( .D(_00895_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5861] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_168 ( .D(_00896_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3716] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1680 ( .D(_00897_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5860] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1681 ( .D(_00898_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5859] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1682 ( .D(_00899_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5858] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1683 ( .D(_00900_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5857] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1684 ( .D(_00901_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5856] ), .QN(_11774_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1685 ( .D(_00902_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5831] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1686 ( .D(_00903_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5830] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1687 ( .D(_00904_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5829] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1688 ( .D(_00905_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5828] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1689 ( .D(_00906_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5827] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_169 ( .D(_00907_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3715] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1690 ( .D(_00908_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5826] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1691 ( .D(_00909_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5825] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1692 ( .D(_00910_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5824] ), .QN(_11773_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1693 ( .D(_00911_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5799] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1694 ( .D(_00912_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5798] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1695 ( .D(_00913_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5797] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1696 ( .D(_00914_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5796] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1697 ( .D(_00915_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5795] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1698 ( .D(_00916_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5794] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1699 ( .D(_00917_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5793] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_17 ( .D(_00918_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4323] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_170 ( .D(_00919_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3714] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1700 ( .D(_00920_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5792] ), .QN(_11772_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1701 ( .D(_00921_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5767] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1702 ( .D(_00922_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5766] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1703 ( .D(_00923_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5765] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1704 ( .D(_00924_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5764] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1705 ( .D(_00925_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5763] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1706 ( .D(_00926_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5762] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1707 ( .D(_00927_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5761] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1708 ( .D(_00928_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5760] ), .QN(_11771_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1709 ( .D(_00929_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5735] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_171 ( .D(_00930_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3713] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1710 ( .D(_00931_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5734] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1711 ( .D(_00932_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5733] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1712 ( .D(_00933_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5732] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1713 ( .D(_00934_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5731] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1714 ( .D(_00935_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5730] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1715 ( .D(_00936_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5729] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1716 ( .D(_00937_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5728] ), .QN(_11770_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1717 ( .D(_00938_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5703] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1718 ( .D(_00939_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5702] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1719 ( .D(_00940_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5701] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_172 ( .D(_00941_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3712] ), .QN(_11769_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1720 ( .D(_00942_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5700] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1721 ( .D(_00943_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5699] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1722 ( .D(_00944_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5698] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1723 ( .D(_00945_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5697] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1724 ( .D(_00946_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5696] ), .QN(_11768_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1725 ( .D(_00947_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5671] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1726 ( .D(_00948_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5670] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1727 ( .D(_00949_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5669] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1728 ( .D(_00950_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5668] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1729 ( .D(_00951_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5667] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_173 ( .D(_00952_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3687] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1730 ( .D(_00953_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5666] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1731 ( .D(_00954_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5665] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1732 ( .D(_00955_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5664] ), .QN(_11767_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1733 ( .D(_00956_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5639] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1734 ( .D(_00957_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5638] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1735 ( .D(_00958_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5637] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1736 ( .D(_00959_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5636] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1737 ( .D(_00960_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5635] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1738 ( .D(_00961_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5634] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1739 ( .D(_00962_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5633] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_174 ( .D(_00963_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3686] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1740 ( .D(_00964_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5632] ), .QN(_11766_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1741 ( .D(_00965_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5607] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1742 ( .D(_00966_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5606] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1743 ( .D(_00967_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5605] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1744 ( .D(_00968_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5604] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1745 ( .D(_00969_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5603] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1746 ( .D(_00970_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5602] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1747 ( .D(_00971_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5601] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1748 ( .D(_00972_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5600] ), .QN(_11765_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1749 ( .D(_00973_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5575] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_175 ( .D(_00974_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3685] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1750 ( .D(_00975_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5574] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1751 ( .D(_00976_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5573] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1752 ( .D(_00977_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5572] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1753 ( .D(_00978_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5571] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1754 ( .D(_00979_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5570] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1755 ( .D(_00980_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5569] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1756 ( .D(_00981_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5568] ), .QN(_11764_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1757 ( .D(_00982_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5543] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1758 ( .D(_00983_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5542] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1759 ( .D(_00984_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5541] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_176 ( .D(_00985_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3684] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1760 ( .D(_00986_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5540] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1761 ( .D(_00987_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5539] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1762 ( .D(_00988_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5538] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1763 ( .D(_00989_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5537] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1764 ( .D(_00990_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5536] ), .QN(_11763_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1765 ( .D(_00991_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5511] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1766 ( .D(_00992_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5510] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1767 ( .D(_00993_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5509] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1768 ( .D(_00994_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5508] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1769 ( .D(_00995_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5507] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_177 ( .D(_00996_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3683] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1770 ( .D(_00997_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5506] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1771 ( .D(_00998_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5505] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1772 ( .D(_00999_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5504] ), .QN(_11762_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1773 ( .D(_01000_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5479] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1774 ( .D(_01001_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5478] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1775 ( .D(_01002_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5477] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1776 ( .D(_01003_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5476] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1777 ( .D(_01004_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5475] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1778 ( .D(_01005_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5474] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1779 ( .D(_01006_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5473] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_178 ( .D(_01007_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3682] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1780 ( .D(_01008_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5472] ), .QN(_11761_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1781 ( .D(_01009_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5447] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1782 ( .D(_01010_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5446] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1783 ( .D(_01011_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5445] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1784 ( .D(_01012_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5444] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1785 ( .D(_01013_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5443] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1786 ( .D(_01014_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5442] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1787 ( .D(_01015_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5441] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1788 ( .D(_01016_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5440] ), .QN(_11760_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1789 ( .D(_01017_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5415] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_179 ( .D(_01018_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3681] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1790 ( .D(_01019_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5414] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1791 ( .D(_01020_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5413] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1792 ( .D(_01021_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5412] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1793 ( .D(_01022_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5411] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1794 ( .D(_01023_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5410] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1795 ( .D(_01024_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5409] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1796 ( .D(_01025_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5408] ), .QN(_11759_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1797 ( .D(_01026_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5383] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1798 ( .D(_01027_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5382] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1799 ( .D(_01028_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5381] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_18 ( .D(_01029_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4322] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_180 ( .D(_01030_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3680] ), .QN(_11758_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1800 ( .D(_01031_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5380] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1801 ( .D(_01032_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5379] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1802 ( .D(_01033_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5378] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1803 ( .D(_01034_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5377] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1804 ( .D(_01035_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5376] ), .QN(_11757_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1805 ( .D(_01036_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5351] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1806 ( .D(_01037_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5350] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1807 ( .D(_01038_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5349] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1808 ( .D(_01039_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5348] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1809 ( .D(_01040_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5347] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_181 ( .D(_01041_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3655] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1810 ( .D(_01042_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5346] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1811 ( .D(_01043_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5345] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1812 ( .D(_01044_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5344] ), .QN(_11756_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1813 ( .D(_01045_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5319] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1814 ( .D(_01046_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5318] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1815 ( .D(_01047_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5317] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1816 ( .D(_01048_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5316] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1817 ( .D(_01049_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5315] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1818 ( .D(_01050_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5314] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1819 ( .D(_01051_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5313] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_182 ( .D(_01052_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3654] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1820 ( .D(_01053_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5312] ), .QN(_11755_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1821 ( .D(_01054_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5287] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1822 ( .D(_01055_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5286] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1823 ( .D(_01056_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5285] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1824 ( .D(_01057_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5284] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1825 ( .D(_01058_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5283] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1826 ( .D(_01059_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5282] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1827 ( .D(_01060_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5281] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1828 ( .D(_01061_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5280] ), .QN(_11754_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1829 ( .D(_01062_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5255] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_183 ( .D(_01063_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3653] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1830 ( .D(_01064_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5254] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1831 ( .D(_01065_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5253] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1832 ( .D(_01066_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5252] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1833 ( .D(_01067_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5251] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1834 ( .D(_01068_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5250] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1835 ( .D(_01069_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5249] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1836 ( .D(_01070_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5248] ), .QN(_11753_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1837 ( .D(_01071_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5223] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1838 ( .D(_01072_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5222] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1839 ( .D(_01073_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5221] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_184 ( .D(_01074_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3652] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1840 ( .D(_01075_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5220] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1841 ( .D(_01076_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5219] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1842 ( .D(_01077_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5218] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1843 ( .D(_01078_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5217] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1844 ( .D(_01079_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5216] ), .QN(_11752_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1845 ( .D(_01080_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5191] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1846 ( .D(_01081_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5190] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1847 ( .D(_01082_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5189] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1848 ( .D(_01083_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5188] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1849 ( .D(_01084_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5187] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_185 ( .D(_01085_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3651] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1850 ( .D(_01086_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5186] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1851 ( .D(_01087_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5185] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1852 ( .D(_01088_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5184] ), .QN(_11751_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1853 ( .D(_01089_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5159] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1854 ( .D(_01090_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5158] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1855 ( .D(_01091_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5157] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1856 ( .D(_01092_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5156] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1857 ( .D(_01093_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5155] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1858 ( .D(_01094_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5154] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1859 ( .D(_01095_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5153] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_186 ( .D(_01096_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3650] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1860 ( .D(_01097_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5152] ), .QN(_11750_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1861 ( .D(_01098_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5127] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1862 ( .D(_01099_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5126] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1863 ( .D(_01100_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5125] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1864 ( .D(_01101_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5124] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1865 ( .D(_01102_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5123] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1866 ( .D(_01103_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5122] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1867 ( .D(_01104_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5121] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1868 ( .D(_01105_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5120] ), .QN(_11749_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1869 ( .D(_01106_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5095] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_187 ( .D(_01107_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3649] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1870 ( .D(_01108_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5094] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1871 ( .D(_01109_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5093] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1872 ( .D(_01110_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5092] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1873 ( .D(_01111_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5091] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1874 ( .D(_01112_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5090] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1875 ( .D(_01113_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5089] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1876 ( .D(_01114_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5088] ), .QN(_11748_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1877 ( .D(_01115_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5063] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1878 ( .D(_01116_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5062] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1879 ( .D(_01117_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5061] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_188 ( .D(_01118_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3648] ), .QN(_11747_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1880 ( .D(_01119_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5060] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1881 ( .D(_01120_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5059] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1882 ( .D(_01121_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5058] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1883 ( .D(_01122_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5057] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1884 ( .D(_01123_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5056] ), .QN(_11746_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1885 ( .D(_01124_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5031] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1886 ( .D(_01125_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5030] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1887 ( .D(_01126_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5029] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1888 ( .D(_01127_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5028] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1889 ( .D(_01128_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5027] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_189 ( .D(_01129_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3623] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1890 ( .D(_01130_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5026] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1891 ( .D(_01131_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5025] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1892 ( .D(_01132_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[5024] ), .QN(_11745_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1893 ( .D(_01133_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4999] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1894 ( .D(_01134_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4998] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1895 ( .D(_01135_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4997] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1896 ( .D(_01136_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4996] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1897 ( .D(_01137_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4995] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1898 ( .D(_01138_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4994] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1899 ( .D(_01139_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4993] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_19 ( .D(_01140_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4321] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_190 ( .D(_01141_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3622] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1900 ( .D(_01142_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4992] ), .QN(_11744_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1901 ( .D(_01143_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4967] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1902 ( .D(_01144_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4966] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1903 ( .D(_01145_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4965] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1904 ( .D(_01146_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4964] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1905 ( .D(_01147_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4963] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1906 ( .D(_01148_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4962] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1907 ( .D(_01149_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4961] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1908 ( .D(_01150_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4960] ), .QN(_11743_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1909 ( .D(_01151_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4935] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_191 ( .D(_01152_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3621] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1910 ( .D(_01153_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4934] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1911 ( .D(_01154_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4933] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1912 ( .D(_01155_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4932] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1913 ( .D(_01156_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4931] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1914 ( .D(_01157_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4930] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1915 ( .D(_01158_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4929] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1916 ( .D(_01159_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4928] ), .QN(_11742_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1917 ( .D(_01160_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4903] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1918 ( .D(_01161_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4902] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1919 ( .D(_01162_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4901] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_192 ( .D(_01163_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3620] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1920 ( .D(_01164_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4900] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1921 ( .D(_01165_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4899] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1922 ( .D(_01166_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4898] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1923 ( .D(_01167_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4897] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1924 ( .D(_01168_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4896] ), .QN(_11741_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1925 ( .D(_01169_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4871] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1926 ( .D(_01170_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4870] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1927 ( .D(_01171_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4869] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1928 ( .D(_01172_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4868] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1929 ( .D(_01173_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4867] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_193 ( .D(_01174_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3619] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1930 ( .D(_01175_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4866] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1931 ( .D(_01176_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4865] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1932 ( .D(_01177_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4864] ), .QN(_11740_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1933 ( .D(_01178_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4839] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1934 ( .D(_01179_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4838] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1935 ( .D(_01180_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4837] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1936 ( .D(_01181_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4836] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1937 ( .D(_01182_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4835] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1938 ( .D(_01183_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4834] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1939 ( .D(_01184_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4833] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_194 ( .D(_01185_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3618] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1940 ( .D(_01186_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4832] ), .QN(_11739_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1941 ( .D(_01187_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4807] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1942 ( .D(_01188_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4806] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1943 ( .D(_01189_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4805] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1944 ( .D(_01190_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4804] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1945 ( .D(_01191_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4803] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1946 ( .D(_01192_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4802] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1947 ( .D(_01193_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4801] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1948 ( .D(_01194_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4800] ), .QN(_11738_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1949 ( .D(_01195_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4775] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_195 ( .D(_01196_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3617] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1950 ( .D(_01197_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4774] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1951 ( .D(_01198_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4773] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1952 ( .D(_01199_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4772] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1953 ( .D(_01200_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4771] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1954 ( .D(_01201_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4770] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1955 ( .D(_01202_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4769] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1956 ( .D(_01203_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4768] ), .QN(_11737_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1957 ( .D(_01204_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4743] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1958 ( .D(_01205_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4742] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1959 ( .D(_01206_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4741] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_196 ( .D(_01207_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3616] ), .QN(_11736_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1960 ( .D(_01208_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4740] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1961 ( .D(_01209_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4739] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1962 ( .D(_01210_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4738] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1963 ( .D(_01211_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4737] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1964 ( .D(_01212_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4736] ), .QN(_11735_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1965 ( .D(_01213_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4711] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1966 ( .D(_01214_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4710] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1967 ( .D(_01215_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4709] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1968 ( .D(_01216_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4708] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1969 ( .D(_01217_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4707] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_197 ( .D(_01218_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3591] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1970 ( .D(_01219_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4706] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1971 ( .D(_01220_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4705] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1972 ( .D(_01221_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4704] ), .QN(_11734_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1973 ( .D(_01222_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4679] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1974 ( .D(_01223_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4678] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1975 ( .D(_01224_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4677] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1976 ( .D(_01225_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4676] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1977 ( .D(_01226_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4675] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1978 ( .D(_01227_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4674] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1979 ( .D(_01228_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4673] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_198 ( .D(_01229_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3590] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1980 ( .D(_01230_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4672] ), .QN(_11733_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1981 ( .D(_01231_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4647] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1982 ( .D(_01232_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4646] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1983 ( .D(_01233_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4645] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1984 ( .D(_01234_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4644] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1985 ( .D(_01235_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4643] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1986 ( .D(_01236_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4642] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1987 ( .D(_01237_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4641] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1988 ( .D(_01238_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4640] ), .QN(_11732_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1989 ( .D(_01239_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4615] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_199 ( .D(_01240_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3589] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1990 ( .D(_01241_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4614] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1991 ( .D(_01242_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4613] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1992 ( .D(_01243_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4612] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1993 ( .D(_01244_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4611] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1994 ( .D(_01245_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4610] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1995 ( .D(_01246_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4609] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1996 ( .D(_01247_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4608] ), .QN(_11731_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1997 ( .D(_01248_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4583] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1998 ( .D(_01249_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4582] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_1999 ( .D(_01250_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4581] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2 ( .D(_01251_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4386] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_20 ( .D(_01252_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4320] ), .QN(_11730_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_200 ( .D(_01253_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3588] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2000 ( .D(_01254_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4580] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2001 ( .D(_01255_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4579] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2002 ( .D(_01256_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4578] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2003 ( .D(_01257_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4577] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2004 ( .D(_01258_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4576] ), .QN(_11729_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2005 ( .D(_01259_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4551] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2006 ( .D(_01260_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4550] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2007 ( .D(_01261_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4549] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2008 ( .D(_01262_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4548] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2009 ( .D(_01263_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4547] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_201 ( .D(_01264_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3587] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2010 ( .D(_01265_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4546] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2011 ( .D(_01266_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4545] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2012 ( .D(_01267_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4544] ), .QN(_11728_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2013 ( .D(_01268_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4519] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2014 ( .D(_01269_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4518] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2015 ( .D(_01270_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4517] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2016 ( .D(_01271_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4516] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2017 ( .D(_01272_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4515] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2018 ( .D(_01273_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4514] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2019 ( .D(_01274_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4513] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_202 ( .D(_01275_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3586] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2020 ( .D(_01276_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4512] ), .QN(_11727_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2021 ( .D(_01277_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4487] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2022 ( .D(_01278_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4486] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2023 ( .D(_01279_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4485] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2024 ( .D(_01280_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4484] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2025 ( .D(_01281_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4483] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2026 ( .D(_01282_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4482] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2027 ( .D(_01283_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4481] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2028 ( .D(_01284_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4480] ), .QN(_11726_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2029 ( .D(_01285_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4455] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_203 ( .D(_01286_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3585] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2030 ( .D(_01287_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4454] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2031 ( .D(_01288_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4453] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2032 ( .D(_01289_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4452] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2033 ( .D(_01290_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4451] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2034 ( .D(_01291_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4450] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2035 ( .D(_01292_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4449] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2036 ( .D(_01293_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4448] ), .QN(_11725_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2037 ( .D(_01294_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4423] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2038 ( .D(_01295_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4422] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2039 ( .D(_01296_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4421] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_204 ( .D(_01297_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3584] ), .QN(_11724_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2040 ( .D(_01298_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4420] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2041 ( .D(_01299_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4419] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2042 ( .D(_01300_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4418] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2043 ( .D(_01301_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4417] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2044 ( .D(_01302_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4416] ), .QN(_11723_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2045 ( .D(_01303_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4391] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2046 ( .D(_01304_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4390] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_2047 ( .D(_01305_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4389] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_205 ( .D(_01306_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3559] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_206 ( .D(_01307_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3558] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_207 ( .D(_01308_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3557] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_208 ( .D(_01309_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3556] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_209 ( .D(_01310_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3555] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_21 ( .D(_01311_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4295] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_210 ( .D(_01312_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3554] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_211 ( .D(_01313_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3553] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_212 ( .D(_01314_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3552] ), .QN(_11722_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_213 ( .D(_01315_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3527] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_214 ( .D(_01316_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3526] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_215 ( .D(_01317_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3525] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_216 ( .D(_01318_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3524] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_217 ( .D(_01319_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3523] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_218 ( .D(_01320_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3522] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_219 ( .D(_01321_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3521] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_22 ( .D(_01322_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4294] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_220 ( .D(_01323_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3520] ), .QN(_11721_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_221 ( .D(_01324_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3495] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_222 ( .D(_01325_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3494] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_223 ( .D(_01326_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3493] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_224 ( .D(_01327_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3492] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_225 ( .D(_01328_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3491] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_226 ( .D(_01329_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3490] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_227 ( .D(_01330_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3489] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_228 ( .D(_01331_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3488] ), .QN(_11720_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_229 ( .D(_01332_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3463] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_23 ( .D(_01333_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4293] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_230 ( .D(_01334_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3462] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_231 ( .D(_01335_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3461] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_232 ( .D(_01336_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3460] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_233 ( .D(_01337_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3459] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_234 ( .D(_01338_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3458] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_235 ( .D(_01339_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3457] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_236 ( .D(_01340_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3456] ), .QN(_11719_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_237 ( .D(_01341_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3431] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_238 ( .D(_01342_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3430] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_239 ( .D(_01343_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3429] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_24 ( .D(_01344_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4292] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_240 ( .D(_01345_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3428] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_241 ( .D(_01346_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3427] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_242 ( .D(_01347_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3426] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_243 ( .D(_01348_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3425] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_244 ( .D(_01349_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3424] ), .QN(_11718_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_245 ( .D(_01350_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3399] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_246 ( .D(_01351_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3398] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_247 ( .D(_01352_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3397] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_248 ( .D(_01353_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3396] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_249 ( .D(_01354_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3395] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_25 ( .D(_01355_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4291] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_250 ( .D(_01356_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3394] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_251 ( .D(_01357_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3393] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_252 ( .D(_01358_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3392] ), .QN(_11717_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_253 ( .D(_01359_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3367] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_254 ( .D(_01360_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3366] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_255 ( .D(_01361_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3365] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_256 ( .D(_01362_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3364] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_257 ( .D(_01363_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3363] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_258 ( .D(_01364_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3362] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_259 ( .D(_01365_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3361] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_26 ( .D(_01366_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4290] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_260 ( .D(_01367_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3360] ), .QN(_11716_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_261 ( .D(_01368_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3335] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_262 ( .D(_01369_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3334] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_263 ( .D(_01370_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3333] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_264 ( .D(_01371_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3332] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_265 ( .D(_01372_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3331] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_266 ( .D(_01373_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3330] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_267 ( .D(_01374_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3329] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_268 ( .D(_01375_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3328] ), .QN(_11715_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_269 ( .D(_01376_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3303] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_27 ( .D(_01377_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4289] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_270 ( .D(_01378_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3302] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_271 ( .D(_01379_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3301] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_272 ( .D(_01380_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3300] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_273 ( .D(_01381_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3299] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_274 ( .D(_01382_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3298] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_275 ( .D(_01383_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3297] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_276 ( .D(_01384_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3296] ), .QN(_11714_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_277 ( .D(_01385_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3271] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_278 ( .D(_01386_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3270] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_279 ( .D(_01387_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3269] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_28 ( .D(_01388_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4288] ), .QN(_11713_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_280 ( .D(_01389_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3268] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_281 ( .D(_01390_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3267] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_282 ( .D(_01391_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3266] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_283 ( .D(_01392_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3265] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_284 ( .D(_01393_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3264] ), .QN(_11712_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_285 ( .D(_01394_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3239] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_286 ( .D(_01395_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3238] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_287 ( .D(_01396_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3237] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_288 ( .D(_01397_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3236] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_289 ( .D(_01398_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3235] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_29 ( .D(_01399_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4263] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_290 ( .D(_01400_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3234] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_291 ( .D(_01401_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3233] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_292 ( .D(_01402_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3232] ), .QN(_11711_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_293 ( .D(_01403_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3207] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_294 ( .D(_01404_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3206] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_295 ( .D(_01405_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3205] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_296 ( .D(_01406_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3204] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_297 ( .D(_01407_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3203] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_298 ( .D(_01408_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3202] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_299 ( .D(_01409_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3201] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_3 ( .D(_01410_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4385] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_30 ( .D(_01411_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4262] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_300 ( .D(_01412_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3200] ), .QN(_11710_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_301 ( .D(_01413_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3175] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_302 ( .D(_01414_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3174] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_303 ( .D(_01415_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3173] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_304 ( .D(_01416_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3172] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_305 ( .D(_01417_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3171] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_306 ( .D(_01418_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3170] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_307 ( .D(_01419_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3169] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_308 ( .D(_01420_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3168] ), .QN(_11709_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_309 ( .D(_01421_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3143] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_31 ( .D(_01422_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4261] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_310 ( .D(_01423_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3142] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_311 ( .D(_01424_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3141] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_312 ( .D(_01425_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3140] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_313 ( .D(_01426_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3139] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_314 ( .D(_01427_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3138] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_315 ( .D(_01428_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3137] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_316 ( .D(_01429_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3136] ), .QN(_11708_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_317 ( .D(_01430_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3111] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_318 ( .D(_01431_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3110] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_319 ( .D(_01432_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3109] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_32 ( .D(_01433_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4260] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_320 ( .D(_01434_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3108] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_321 ( .D(_01435_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3107] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_322 ( .D(_01436_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3106] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_323 ( .D(_01437_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3105] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_324 ( .D(_01438_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3104] ), .QN(_11707_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_325 ( .D(_01439_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3079] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_326 ( .D(_01440_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3078] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_327 ( .D(_01441_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3077] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_328 ( .D(_01442_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3076] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_329 ( .D(_01443_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3075] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_33 ( .D(_01444_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4259] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_330 ( .D(_01445_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3074] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_331 ( .D(_01446_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3073] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_332 ( .D(_01447_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3072] ), .QN(_11706_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_333 ( .D(_01448_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3047] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_334 ( .D(_01449_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3046] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_335 ( .D(_01450_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3045] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_336 ( .D(_01451_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3044] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_337 ( .D(_01452_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3043] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_338 ( .D(_01453_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3042] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_339 ( .D(_01454_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3041] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_34 ( .D(_01455_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4258] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_340 ( .D(_01456_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3040] ), .QN(_11705_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_341 ( .D(_01457_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3015] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_342 ( .D(_01458_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3014] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_343 ( .D(_01459_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3013] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_344 ( .D(_01460_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3012] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_345 ( .D(_01461_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3011] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_346 ( .D(_01462_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3010] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_347 ( .D(_01463_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3009] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_348 ( .D(_01464_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[3008] ), .QN(_11704_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_349 ( .D(_01465_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2983] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_35 ( .D(_01466_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4257] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_350 ( .D(_01467_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2982] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_351 ( .D(_01468_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2981] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_352 ( .D(_01469_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2980] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_353 ( .D(_01470_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2979] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_354 ( .D(_01471_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2978] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_355 ( .D(_01472_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2977] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_356 ( .D(_01473_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2976] ), .QN(_11703_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_357 ( .D(_01474_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2951] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_358 ( .D(_01475_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2950] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_359 ( .D(_01476_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2949] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_36 ( .D(_01477_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4256] ), .QN(_11702_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_360 ( .D(_01478_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2948] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_361 ( .D(_01479_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2947] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_362 ( .D(_01480_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2946] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_363 ( .D(_01481_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2945] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_364 ( .D(_01482_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2944] ), .QN(_11701_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_365 ( .D(_01483_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2919] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_366 ( .D(_01484_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2918] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_367 ( .D(_01485_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2917] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_368 ( .D(_01486_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2916] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_369 ( .D(_01487_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2915] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_37 ( .D(_01488_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4231] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_370 ( .D(_01489_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2914] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_371 ( .D(_01490_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2913] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_372 ( .D(_01491_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2912] ), .QN(_11700_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_373 ( .D(_01492_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2887] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_374 ( .D(_01493_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2886] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_375 ( .D(_01494_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2885] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_376 ( .D(_01495_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2884] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_377 ( .D(_01496_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2883] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_378 ( .D(_01497_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2882] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_379 ( .D(_01498_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2881] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_38 ( .D(_01499_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4230] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_380 ( .D(_01500_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2880] ), .QN(_11699_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_381 ( .D(_01501_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2855] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_382 ( .D(_01502_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2854] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_383 ( .D(_01503_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2853] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_384 ( .D(_01504_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2852] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_385 ( .D(_01505_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2851] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_386 ( .D(_01506_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2850] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_387 ( .D(_01507_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2849] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_388 ( .D(_01508_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2848] ), .QN(_11698_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_389 ( .D(_01509_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2823] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_39 ( .D(_01510_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4229] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_390 ( .D(_01511_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2822] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_391 ( .D(_01512_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2821] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_392 ( .D(_01513_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2820] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_393 ( .D(_01514_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2819] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_394 ( .D(_01515_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2818] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_395 ( .D(_01516_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2817] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_396 ( .D(_01517_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2816] ), .QN(_11697_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_397 ( .D(_01518_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2791] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_398 ( .D(_01519_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2790] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_399 ( .D(_01520_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2789] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_4 ( .D(_01521_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4384] ), .QN(_11696_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_40 ( .D(_01522_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4228] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_400 ( .D(_01523_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2788] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_401 ( .D(_01524_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2787] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_402 ( .D(_01525_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2786] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_403 ( .D(_01526_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2785] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_404 ( .D(_01527_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2784] ), .QN(_11695_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_405 ( .D(_01528_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2759] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_406 ( .D(_01529_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2758] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_407 ( .D(_01530_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2757] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_408 ( .D(_01531_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2756] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_409 ( .D(_01532_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2755] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_41 ( .D(_01533_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4227] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_410 ( .D(_01534_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2754] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_411 ( .D(_01535_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2753] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_412 ( .D(_01536_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2752] ), .QN(_11694_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_413 ( .D(_01537_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2727] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_414 ( .D(_01538_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2726] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_415 ( .D(_01539_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2725] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_416 ( .D(_01540_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2724] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_417 ( .D(_01541_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2723] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_418 ( .D(_01542_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2722] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_419 ( .D(_01543_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2721] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_42 ( .D(_01544_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4226] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_420 ( .D(_01545_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2720] ), .QN(_11693_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_421 ( .D(_01546_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2695] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_422 ( .D(_01547_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2694] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_423 ( .D(_01548_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2693] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_424 ( .D(_01549_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2692] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_425 ( .D(_01550_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2691] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_426 ( .D(_01551_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2690] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_427 ( .D(_01552_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2689] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_428 ( .D(_01553_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2688] ), .QN(_11692_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_429 ( .D(_01554_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2663] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_43 ( .D(_01555_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4225] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_430 ( .D(_01556_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2662] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_431 ( .D(_01557_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2661] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_432 ( .D(_01558_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2660] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_433 ( .D(_01559_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2659] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_434 ( .D(_01560_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2658] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_435 ( .D(_01561_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2657] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_436 ( .D(_01562_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2656] ), .QN(_11691_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_437 ( .D(_01563_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2631] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_438 ( .D(_01564_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2630] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_439 ( .D(_01565_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2629] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_44 ( .D(_01566_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4224] ), .QN(_11690_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_440 ( .D(_01567_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2628] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_441 ( .D(_01568_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2627] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_442 ( .D(_01569_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2626] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_443 ( .D(_01570_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2625] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_444 ( .D(_01571_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2624] ), .QN(_11689_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_445 ( .D(_01572_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2599] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_446 ( .D(_01573_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2598] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_447 ( .D(_01574_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2597] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_448 ( .D(_01575_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2596] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_449 ( .D(_01576_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2595] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_45 ( .D(_01577_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4199] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_450 ( .D(_01578_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2594] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_451 ( .D(_01579_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2593] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_452 ( .D(_01580_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2592] ), .QN(_11688_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_453 ( .D(_01581_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2567] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_454 ( .D(_01582_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2566] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_455 ( .D(_01583_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2565] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_456 ( .D(_01584_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2564] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_457 ( .D(_01585_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2563] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_458 ( .D(_01586_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2562] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_459 ( .D(_01587_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2561] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_46 ( .D(_01588_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4198] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_460 ( .D(_01589_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2560] ), .QN(_11687_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_461 ( .D(_01590_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2535] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_462 ( .D(_01591_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2534] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_463 ( .D(_01592_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2533] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_464 ( .D(_01593_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2532] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_465 ( .D(_01594_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2531] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_466 ( .D(_01595_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2530] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_467 ( .D(_01596_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2529] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_468 ( .D(_01597_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2528] ), .QN(_11686_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_469 ( .D(_01598_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2503] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_47 ( .D(_01599_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4197] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_470 ( .D(_01600_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2502] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_471 ( .D(_01601_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2501] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_472 ( .D(_01602_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2500] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_473 ( .D(_01603_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2499] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_474 ( .D(_01604_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2498] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_475 ( .D(_01605_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2497] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_476 ( .D(_01606_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2496] ), .QN(_11685_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_477 ( .D(_01607_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2471] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_478 ( .D(_01608_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2470] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_479 ( .D(_01609_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2469] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_48 ( .D(_01610_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4196] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_480 ( .D(_01611_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2468] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_481 ( .D(_01612_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2467] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_482 ( .D(_01613_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2466] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_483 ( .D(_01614_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2465] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_484 ( .D(_01615_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2464] ), .QN(_11684_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_485 ( .D(_01616_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2439] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_486 ( .D(_01617_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2438] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_487 ( .D(_01618_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2437] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_488 ( .D(_01619_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2436] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_489 ( .D(_01620_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2435] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_49 ( .D(_01621_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4195] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_490 ( .D(_01622_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2434] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_491 ( .D(_01623_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2433] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_492 ( .D(_01624_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2432] ), .QN(_11683_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_493 ( .D(_01625_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2407] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_494 ( .D(_01626_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2406] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_495 ( .D(_01627_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2405] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_496 ( .D(_01628_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2404] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_497 ( .D(_01629_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2403] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_498 ( .D(_01630_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2402] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_499 ( .D(_01631_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2401] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_5 ( .D(_01632_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4359] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_50 ( .D(_01633_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4194] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_500 ( .D(_01634_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2400] ), .QN(_11682_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_501 ( .D(_01635_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2375] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_502 ( .D(_01636_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2374] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_503 ( .D(_01637_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2373] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_504 ( .D(_01638_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2372] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_505 ( .D(_01639_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2371] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_506 ( .D(_01640_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2370] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_507 ( .D(_01641_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2369] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_508 ( .D(_01642_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2368] ), .QN(_11681_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_509 ( .D(_01643_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2343] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_51 ( .D(_01644_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4193] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_510 ( .D(_01645_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2342] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_511 ( .D(_01646_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2341] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_512 ( .D(_01647_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2340] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_513 ( .D(_01648_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2339] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_514 ( .D(_01649_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2338] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_515 ( .D(_01650_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2337] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_516 ( .D(_01651_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2336] ), .QN(_11680_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_517 ( .D(_01652_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2311] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_518 ( .D(_01653_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2310] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_519 ( .D(_01654_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2309] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_52 ( .D(_01655_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4192] ), .QN(_11679_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_520 ( .D(_01656_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2308] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_521 ( .D(_01657_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2307] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_522 ( .D(_01658_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2306] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_523 ( .D(_01659_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2305] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_524 ( .D(_01660_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2304] ), .QN(_11678_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_525 ( .D(_01661_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2279] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_526 ( .D(_01662_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2278] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_527 ( .D(_01663_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2277] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_528 ( .D(_01664_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2276] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_529 ( .D(_01665_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2275] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_53 ( .D(_01666_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4167] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_530 ( .D(_01667_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2274] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_531 ( .D(_01668_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2273] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_532 ( .D(_01669_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2272] ), .QN(_11677_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_533 ( .D(_01670_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2247] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_534 ( .D(_01671_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2246] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_535 ( .D(_01672_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2245] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_536 ( .D(_01673_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2244] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_537 ( .D(_01674_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2243] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_538 ( .D(_01675_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2242] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_539 ( .D(_01676_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2241] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_54 ( .D(_01677_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4166] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_540 ( .D(_01678_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2240] ), .QN(_11676_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_541 ( .D(_01679_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2215] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_542 ( .D(_01680_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2214] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_543 ( .D(_01681_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2213] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_544 ( .D(_01682_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2212] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_545 ( .D(_01683_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2211] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_546 ( .D(_01684_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2210] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_547 ( .D(_01685_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2209] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_548 ( .D(_01686_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2208] ), .QN(_11675_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_549 ( .D(_01687_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2183] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_55 ( .D(_01688_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4165] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_550 ( .D(_01689_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2182] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_551 ( .D(_01690_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2181] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_552 ( .D(_01691_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2180] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_553 ( .D(_01692_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2179] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_554 ( .D(_01693_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2178] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_555 ( .D(_01694_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2177] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_556 ( .D(_01695_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2176] ), .QN(_11674_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_557 ( .D(_01696_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2151] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_558 ( .D(_01697_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2150] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_559 ( .D(_01698_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2149] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_56 ( .D(_01699_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4164] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_560 ( .D(_01700_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2148] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_561 ( .D(_01701_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2147] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_562 ( .D(_01702_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2146] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_563 ( .D(_01703_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2145] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_564 ( .D(_01704_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2144] ), .QN(_11673_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_565 ( .D(_01705_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2119] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_566 ( .D(_01706_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2118] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_567 ( .D(_01707_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2117] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_568 ( .D(_01708_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2116] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_569 ( .D(_01709_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2115] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_57 ( .D(_01710_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4163] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_570 ( .D(_01711_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2114] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_571 ( .D(_01712_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2113] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_572 ( .D(_01713_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2112] ), .QN(_11672_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_573 ( .D(_01714_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2087] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_574 ( .D(_01715_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2086] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_575 ( .D(_01716_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2085] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_576 ( .D(_01717_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2084] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_577 ( .D(_01718_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2083] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_578 ( .D(_01719_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2082] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_579 ( .D(_01720_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2081] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_58 ( .D(_01721_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4162] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_580 ( .D(_01722_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2080] ), .QN(_11671_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_581 ( .D(_01723_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2055] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_582 ( .D(_01724_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2054] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_583 ( .D(_01725_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2053] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_584 ( .D(_01726_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2052] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_585 ( .D(_01727_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2051] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_586 ( .D(_01728_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2050] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_587 ( .D(_01729_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2049] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_588 ( .D(_01730_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2048] ), .QN(_11670_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_589 ( .D(_01731_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2023] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_59 ( .D(_01732_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4161] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_590 ( .D(_01733_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2022] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_591 ( .D(_01734_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2021] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_592 ( .D(_01735_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2020] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_593 ( .D(_01736_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2019] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_594 ( .D(_01737_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2018] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_595 ( .D(_01738_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2017] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_596 ( .D(_01739_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[2016] ), .QN(_11669_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_597 ( .D(_01740_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1991] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_598 ( .D(_01741_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1990] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_599 ( .D(_01742_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1989] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_6 ( .D(_01743_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4358] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_60 ( .D(_01744_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4160] ), .QN(_11668_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_600 ( .D(_01745_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1988] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_601 ( .D(_01746_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1987] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_602 ( .D(_01747_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1986] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_603 ( .D(_01748_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1985] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_604 ( .D(_01749_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1984] ), .QN(_11667_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_605 ( .D(_01750_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1959] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_606 ( .D(_01751_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1958] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_607 ( .D(_01752_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1957] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_608 ( .D(_01753_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1956] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_609 ( .D(_01754_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1955] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_61 ( .D(_01755_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4135] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_610 ( .D(_01756_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1954] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_611 ( .D(_01757_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1953] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_612 ( .D(_01758_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1952] ), .QN(_11666_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_613 ( .D(_01759_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1927] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_614 ( .D(_01760_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1926] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_615 ( .D(_01761_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1925] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_616 ( .D(_01762_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1924] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_617 ( .D(_01763_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1923] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_618 ( .D(_01764_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1922] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_619 ( .D(_01765_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1921] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_62 ( .D(_01766_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4134] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_620 ( .D(_01767_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1920] ), .QN(_11665_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_621 ( .D(_01768_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1895] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_622 ( .D(_01769_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1894] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_623 ( .D(_01770_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1893] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_624 ( .D(_01771_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1892] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_625 ( .D(_01772_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1891] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_626 ( .D(_01773_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1890] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_627 ( .D(_01774_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1889] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_628 ( .D(_01775_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1888] ), .QN(_11664_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_629 ( .D(_01776_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1863] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_63 ( .D(_01777_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4133] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_630 ( .D(_01778_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1862] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_631 ( .D(_01779_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1861] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_632 ( .D(_01780_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1860] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_633 ( .D(_01781_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1859] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_634 ( .D(_01782_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1858] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_635 ( .D(_01783_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1857] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_636 ( .D(_01784_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1856] ), .QN(_11663_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_637 ( .D(_01785_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1831] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_638 ( .D(_01786_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1830] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_639 ( .D(_01787_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1829] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_64 ( .D(_01788_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4132] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_640 ( .D(_01789_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1828] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_641 ( .D(_01790_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1827] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_642 ( .D(_01791_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1826] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_643 ( .D(_01792_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1825] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_644 ( .D(_01793_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1824] ), .QN(_11662_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_645 ( .D(_01794_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1799] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_646 ( .D(_01795_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1798] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_647 ( .D(_01796_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1797] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_648 ( .D(_01797_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1796] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_649 ( .D(_01798_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1795] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_65 ( .D(_01799_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4131] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_650 ( .D(_01800_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1794] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_651 ( .D(_01801_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1793] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_652 ( .D(_01802_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1792] ), .QN(_11661_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_653 ( .D(_01803_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1767] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_654 ( .D(_01804_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1766] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_655 ( .D(_01805_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1765] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_656 ( .D(_01806_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1764] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_657 ( .D(_01807_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1763] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_658 ( .D(_01808_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1762] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_659 ( .D(_01809_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1761] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_66 ( .D(_01810_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4130] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_660 ( .D(_01811_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1760] ), .QN(_11660_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_661 ( .D(_01812_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1735] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_662 ( .D(_01813_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1734] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_663 ( .D(_01814_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1733] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_664 ( .D(_01815_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1732] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_665 ( .D(_01816_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1731] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_666 ( .D(_01817_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1730] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_667 ( .D(_01818_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1729] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_668 ( .D(_01819_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1728] ), .QN(_11659_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_669 ( .D(_01820_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1703] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_67 ( .D(_01821_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4129] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_670 ( .D(_01822_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1702] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_671 ( .D(_01823_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1701] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_672 ( .D(_01824_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1700] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_673 ( .D(_01825_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1699] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_674 ( .D(_01826_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1698] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_675 ( .D(_01827_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1697] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_676 ( .D(_01828_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1696] ), .QN(_11658_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_677 ( .D(_01829_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1671] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_678 ( .D(_01830_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1670] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_679 ( .D(_01831_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1669] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_68 ( .D(_01832_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4128] ), .QN(_11657_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_680 ( .D(_01833_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1668] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_681 ( .D(_01834_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1667] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_682 ( .D(_01835_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1666] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_683 ( .D(_01836_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1665] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_684 ( .D(_01837_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1664] ), .QN(_11656_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_685 ( .D(_01838_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1639] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_686 ( .D(_01839_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1638] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_687 ( .D(_01840_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1637] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_688 ( .D(_01841_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1636] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_689 ( .D(_01842_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1635] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_69 ( .D(_01843_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4103] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_690 ( .D(_01844_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1634] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_691 ( .D(_01845_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1633] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_692 ( .D(_01846_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1632] ), .QN(_11655_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_693 ( .D(_01847_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1607] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_694 ( .D(_01848_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1606] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_695 ( .D(_01849_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1605] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_696 ( .D(_01850_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1604] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_697 ( .D(_01851_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1603] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_698 ( .D(_01852_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1602] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_699 ( .D(_01853_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1601] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_7 ( .D(_01854_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4357] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_70 ( .D(_01855_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4102] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_700 ( .D(_01856_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1600] ), .QN(_11654_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_701 ( .D(_01857_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1575] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_702 ( .D(_01858_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1574] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_703 ( .D(_01859_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1573] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_704 ( .D(_01860_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1572] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_705 ( .D(_01861_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1571] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_706 ( .D(_01862_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1570] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_707 ( .D(_01863_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1569] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_708 ( .D(_01864_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1568] ), .QN(_11653_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_709 ( .D(_01865_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1543] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_71 ( .D(_01866_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4101] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_710 ( .D(_01867_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1542] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_711 ( .D(_01868_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1541] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_712 ( .D(_01869_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1540] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_713 ( .D(_01870_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1539] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_714 ( .D(_01871_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1538] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_715 ( .D(_01872_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1537] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_716 ( .D(_01873_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1536] ), .QN(_11652_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_717 ( .D(_01874_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1511] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_718 ( .D(_01875_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1510] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_719 ( .D(_01876_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1509] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_72 ( .D(_01877_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4100] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_720 ( .D(_01878_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1508] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_721 ( .D(_01879_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1507] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_722 ( .D(_01880_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1506] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_723 ( .D(_01881_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1505] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_724 ( .D(_01882_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1504] ), .QN(_11651_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_725 ( .D(_01883_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1479] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_726 ( .D(_01884_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1478] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_727 ( .D(_01885_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1477] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_728 ( .D(_01886_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1476] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_729 ( .D(_01887_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1475] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_73 ( .D(_01888_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4099] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_730 ( .D(_01889_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1474] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_731 ( .D(_01890_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1473] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_732 ( .D(_01891_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1472] ), .QN(_11650_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_733 ( .D(_01892_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1447] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_734 ( .D(_01893_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1446] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_735 ( .D(_01894_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1445] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_736 ( .D(_01895_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1444] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_737 ( .D(_01896_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1443] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_738 ( .D(_01897_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1442] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_739 ( .D(_01898_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1441] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_74 ( .D(_01899_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4098] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_740 ( .D(_01900_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1440] ), .QN(_11649_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_741 ( .D(_01901_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1415] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_742 ( .D(_01902_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1414] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_743 ( .D(_01903_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1413] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_744 ( .D(_01904_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1412] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_745 ( .D(_01905_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1411] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_746 ( .D(_01906_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1410] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_747 ( .D(_01907_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1409] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_748 ( .D(_01908_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1408] ), .QN(_11648_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_749 ( .D(_01909_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1383] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_75 ( .D(_01910_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4097] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_750 ( .D(_01911_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1382] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_751 ( .D(_01912_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1381] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_752 ( .D(_01913_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1380] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_753 ( .D(_01914_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1379] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_754 ( .D(_01915_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1378] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_755 ( .D(_01916_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1377] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_756 ( .D(_01917_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1376] ), .QN(_11647_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_757 ( .D(_01918_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1351] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_758 ( .D(_01919_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1350] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_759 ( .D(_01920_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1349] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_76 ( .D(_01921_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4096] ), .QN(_11646_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_760 ( .D(_01922_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1348] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_761 ( .D(_01923_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1347] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_762 ( .D(_01924_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1346] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_763 ( .D(_01925_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1345] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_764 ( .D(_01926_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1344] ), .QN(_11645_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_765 ( .D(_01927_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1319] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_766 ( .D(_01928_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1318] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_767 ( .D(_01929_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1317] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_768 ( .D(_01930_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1316] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_769 ( .D(_01931_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1315] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_77 ( .D(_01932_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4071] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_770 ( .D(_01933_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1314] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_771 ( .D(_01934_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1313] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_772 ( .D(_01935_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1312] ), .QN(_11644_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_773 ( .D(_01936_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1287] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_774 ( .D(_01937_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1286] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_775 ( .D(_01938_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1285] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_776 ( .D(_01939_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1284] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_777 ( .D(_01940_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1283] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_778 ( .D(_01941_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1282] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_779 ( .D(_01942_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1281] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_78 ( .D(_01943_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4070] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_780 ( .D(_01944_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1280] ), .QN(_11643_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_781 ( .D(_01945_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1255] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_782 ( .D(_01946_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1254] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_783 ( .D(_01947_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1253] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_784 ( .D(_01948_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1252] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_785 ( .D(_01949_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1251] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_786 ( .D(_01950_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1250] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_787 ( .D(_01951_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1249] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_788 ( .D(_01952_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1248] ), .QN(_11642_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_789 ( .D(_01953_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1223] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_79 ( .D(_01954_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4069] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_790 ( .D(_01955_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1222] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_791 ( .D(_01956_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1221] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_792 ( .D(_01957_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1220] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_793 ( .D(_01958_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1219] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_794 ( .D(_01959_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1218] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_795 ( .D(_01960_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1217] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_796 ( .D(_01961_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1216] ), .QN(_11641_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_797 ( .D(_01962_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1191] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_798 ( .D(_01963_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1190] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_799 ( .D(_01964_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1189] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_8 ( .D(_01965_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4356] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_80 ( .D(_01966_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4068] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_800 ( .D(_01967_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1188] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_801 ( .D(_01968_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1187] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_802 ( .D(_01969_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1186] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_803 ( .D(_01970_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1185] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_804 ( .D(_01971_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1184] ), .QN(_11640_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_805 ( .D(_01972_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1159] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_806 ( .D(_01973_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1158] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_807 ( .D(_01974_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1157] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_808 ( .D(_01975_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1156] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_809 ( .D(_01976_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1155] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_81 ( .D(_01977_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4067] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_810 ( .D(_01978_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1154] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_811 ( .D(_01979_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1153] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_812 ( .D(_01980_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1152] ), .QN(_11639_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_813 ( .D(_01981_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1127] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_814 ( .D(_01982_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1126] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_815 ( .D(_01983_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1125] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_816 ( .D(_01984_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1124] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_817 ( .D(_01985_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1123] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_818 ( .D(_01986_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1122] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_819 ( .D(_01987_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1121] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_82 ( .D(_01988_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4066] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_820 ( .D(_01989_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1120] ), .QN(_11638_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_821 ( .D(_01990_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1095] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_822 ( .D(_01991_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1094] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_823 ( .D(_01992_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1093] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_824 ( .D(_01993_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1092] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_825 ( .D(_01994_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1091] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_826 ( .D(_01995_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1090] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_827 ( .D(_01996_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1089] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_828 ( .D(_01997_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1088] ), .QN(_11637_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_829 ( .D(_01998_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1063] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_83 ( .D(_01999_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4065] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_830 ( .D(_02000_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1062] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_831 ( .D(_02001_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1061] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_832 ( .D(_02002_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1060] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_833 ( .D(_02003_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1059] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_834 ( .D(_02004_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1058] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_835 ( .D(_02005_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1057] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_836 ( .D(_02006_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1056] ), .QN(_11636_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_837 ( .D(_02007_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1031] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_838 ( .D(_02008_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1030] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_839 ( .D(_02009_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1029] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_84 ( .D(_02010_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4064] ), .QN(_11635_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_840 ( .D(_02011_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1028] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_841 ( .D(_02012_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1027] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_842 ( .D(_02013_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1026] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_843 ( .D(_02014_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1025] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_844 ( .D(_02015_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[1024] ), .QN(_11634_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_845 ( .D(_02016_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[999] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_846 ( .D(_02017_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[998] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_847 ( .D(_02018_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[997] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_848 ( .D(_02019_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[996] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_849 ( .D(_02020_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[995] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_85 ( .D(_02021_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4039] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_850 ( .D(_02022_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[994] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_851 ( .D(_02023_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[993] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_852 ( .D(_02024_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[992] ), .QN(_11633_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_853 ( .D(_02025_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[967] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_854 ( .D(_02026_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[966] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_855 ( .D(_02027_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[965] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_856 ( .D(_02028_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[964] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_857 ( .D(_02029_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[963] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_858 ( .D(_02030_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[962] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_859 ( .D(_02031_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[961] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_86 ( .D(_02032_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4038] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_860 ( .D(_02033_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[960] ), .QN(_11632_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_861 ( .D(_02034_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[935] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_862 ( .D(_02035_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[934] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_863 ( .D(_02036_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[933] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_864 ( .D(_02037_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[932] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_865 ( .D(_02038_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[931] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_866 ( .D(_02039_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[930] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_867 ( .D(_02040_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[929] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_868 ( .D(_02041_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[928] ), .QN(_11631_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_869 ( .D(_02042_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[903] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_87 ( .D(_02043_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4037] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_870 ( .D(_02044_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[902] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_871 ( .D(_02045_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[901] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_872 ( .D(_02046_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[900] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_873 ( .D(_02047_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[899] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_874 ( .D(_02048_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[898] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_875 ( .D(_02049_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[897] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_876 ( .D(_02050_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[896] ), .QN(_11630_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_877 ( .D(_02051_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[871] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_878 ( .D(_02052_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[870] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_879 ( .D(_02053_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[869] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_88 ( .D(_02054_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4036] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_880 ( .D(_02055_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[868] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_881 ( .D(_02056_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[867] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_882 ( .D(_02057_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[866] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_883 ( .D(_02058_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[865] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_884 ( .D(_02059_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[864] ), .QN(_11629_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_885 ( .D(_02060_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[839] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_886 ( .D(_02061_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[838] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_887 ( .D(_02062_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[837] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_888 ( .D(_02063_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[836] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_889 ( .D(_02064_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[835] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_89 ( .D(_02065_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4035] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_890 ( .D(_02066_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[834] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_891 ( .D(_02067_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[833] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_892 ( .D(_02068_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[832] ), .QN(_11628_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_893 ( .D(_02069_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[807] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_894 ( .D(_02070_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[806] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_895 ( .D(_02071_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[805] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_896 ( .D(_02072_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[804] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_897 ( .D(_02073_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[803] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_898 ( .D(_02074_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[802] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_899 ( .D(_02075_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[801] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_9 ( .D(_02076_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4355] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_90 ( .D(_02077_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4034] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_900 ( .D(_02078_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[800] ), .QN(_11627_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_901 ( .D(_02079_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[775] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_902 ( .D(_02080_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[774] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_903 ( .D(_02081_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[773] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_904 ( .D(_02082_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[772] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_905 ( .D(_02083_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[771] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_906 ( .D(_02084_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[770] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_907 ( .D(_02085_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[769] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_908 ( .D(_02086_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[768] ), .QN(_11626_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_909 ( .D(_02087_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[743] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_91 ( .D(_02088_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4033] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_910 ( .D(_02089_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[742] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_911 ( .D(_02090_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[741] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_912 ( .D(_02091_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[740] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_913 ( .D(_02092_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[739] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_914 ( .D(_02093_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[738] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_915 ( .D(_02094_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[737] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_916 ( .D(_02095_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[736] ), .QN(_11625_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_917 ( .D(_02096_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[711] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_918 ( .D(_02097_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[710] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_919 ( .D(_02098_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[709] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_92 ( .D(_02099_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4032] ), .QN(_11624_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_920 ( .D(_02100_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[708] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_921 ( .D(_02101_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[707] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_922 ( .D(_02102_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[706] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_923 ( .D(_02103_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[705] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_924 ( .D(_02104_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[704] ), .QN(_11623_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_925 ( .D(_02105_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[679] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_926 ( .D(_02106_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[678] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_927 ( .D(_02107_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[677] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_928 ( .D(_02108_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[676] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_929 ( .D(_02109_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[675] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_93 ( .D(_02110_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4007] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_930 ( .D(_02111_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[674] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_931 ( .D(_02112_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[673] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_932 ( .D(_02113_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[672] ), .QN(_11622_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_933 ( .D(_02114_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[647] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_934 ( .D(_02115_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[646] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_935 ( .D(_02116_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[645] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_936 ( .D(_02117_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[644] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_937 ( .D(_02118_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[643] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_938 ( .D(_02119_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[642] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_939 ( .D(_02120_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[641] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_94 ( .D(_02121_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4006] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_940 ( .D(_02122_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[640] ), .QN(_11621_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_941 ( .D(_02123_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[615] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_942 ( .D(_02124_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[614] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_943 ( .D(_02125_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[613] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_944 ( .D(_02126_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[612] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_945 ( .D(_02127_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[611] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_946 ( .D(_02128_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[610] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_947 ( .D(_02129_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[609] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_948 ( .D(_02130_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[608] ), .QN(_11620_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_949 ( .D(_02131_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[583] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_95 ( .D(_02132_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4005] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_950 ( .D(_02133_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[582] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_951 ( .D(_02134_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[581] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_952 ( .D(_02135_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[580] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_953 ( .D(_02136_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[579] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_954 ( .D(_02137_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[578] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_955 ( .D(_02138_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[577] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_956 ( .D(_02139_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[576] ), .QN(_11619_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_957 ( .D(_02140_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[551] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_958 ( .D(_02141_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[550] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_959 ( .D(_02142_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[549] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_96 ( .D(_02143_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4004] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_960 ( .D(_02144_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[548] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_961 ( .D(_02145_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[547] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_962 ( .D(_02146_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[546] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_963 ( .D(_02147_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[545] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_964 ( .D(_02148_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[544] ), .QN(_11618_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_965 ( .D(_02149_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[519] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_966 ( .D(_02150_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[518] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_967 ( .D(_02151_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[517] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_968 ( .D(_02152_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[516] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_969 ( .D(_02153_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[515] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_97 ( .D(_02154_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4003] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_970 ( .D(_02155_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[514] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_971 ( .D(_02156_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[513] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_972 ( .D(_02157_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[512] ), .QN(_11617_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_973 ( .D(_02158_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[487] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_974 ( .D(_02159_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[486] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_975 ( .D(_02160_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[485] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_976 ( .D(_02161_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[484] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_977 ( .D(_02162_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[483] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_978 ( .D(_02163_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[482] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_979 ( .D(_02164_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[481] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_98 ( .D(_02165_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4002] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_980 ( .D(_02166_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[480] ), .QN(_11616_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_981 ( .D(_02167_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[455] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_982 ( .D(_02168_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[454] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_983 ( .D(_02169_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[453] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_984 ( .D(_02170_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[452] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_985 ( .D(_02171_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[451] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_986 ( .D(_02172_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[450] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_987 ( .D(_02173_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[449] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_988 ( .D(_02174_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[448] ), .QN(_11615_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_989 ( .D(_02175_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[423] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_99 ( .D(_02176_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[4001] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_990 ( .D(_02177_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[422] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_991 ( .D(_02178_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[421] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_992 ( .D(_02179_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[420] ), .QN(load_data_out_$_NOR__Y_3_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_993 ( .D(_02180_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[419] ), .QN(load_data_out_$_NOR__Y_4_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_994 ( .D(_02181_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[418] ), .QN(load_data_out_$_NOR__Y_5_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_995 ( .D(_02182_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[417] ), .QN(load_data_out_$_NOR__Y_6_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_996 ( .D(_02183_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[416] ), .QN(_11614_ ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_997 ( .D(_02184_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[391] ), .QN(load_data_out_$_NOR__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_998 ( .D(_02185_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[390] ), .QN(load_data_out_$_NOR__Y_1_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \u_lsu.pmem_$_SDFFE_PP0P__Q_999 ( .D(_02186_ ), .CK(_11608_ ), .Q(\u_lsu.pmem[389] ), .QN(load_data_out_$_NOR__Y_2_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
BUF_X8 fanout_buf_1 ( .A(_00000_ ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(\ifu_rdata[15] ), .Z(fanout_net_2 ) );
BUF_X8 fanout_buf_3 ( .A(\ifu_rdata[15] ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(\ifu_rdata[16] ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(\ifu_rdata[20] ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(\ifu_rdata[20] ), .Z(fanout_net_6 ) );
BUF_X8 fanout_buf_7 ( .A(\ifu_rdata[21] ), .Z(fanout_net_7 ) );
BUF_X8 fanout_buf_8 ( .A(fanout_net_75 ), .Z(fanout_net_8 ) );
BUF_X8 fanout_buf_9 ( .A(fanout_net_75 ), .Z(fanout_net_9 ) );
BUF_X8 fanout_buf_10 ( .A(fanout_net_75 ), .Z(fanout_net_10 ) );
BUF_X8 fanout_buf_11 ( .A(fanout_net_75 ), .Z(fanout_net_11 ) );
BUF_X8 fanout_buf_12 ( .A(fanout_net_75 ), .Z(fanout_net_12 ) );
BUF_X8 fanout_buf_13 ( .A(fanout_net_75 ), .Z(fanout_net_13 ) );
BUF_X8 fanout_buf_14 ( .A(fanout_net_75 ), .Z(fanout_net_14 ) );
BUF_X8 fanout_buf_15 ( .A(fanout_net_75 ), .Z(fanout_net_15 ) );
BUF_X8 fanout_buf_16 ( .A(fanout_net_75 ), .Z(fanout_net_16 ) );
BUF_X8 fanout_buf_17 ( .A(fanout_net_75 ), .Z(fanout_net_17 ) );
BUF_X8 fanout_buf_18 ( .A(fanout_net_75 ), .Z(fanout_net_18 ) );
BUF_X8 fanout_buf_19 ( .A(fanout_net_75 ), .Z(fanout_net_19 ) );
BUF_X8 fanout_buf_20 ( .A(fanout_net_75 ), .Z(fanout_net_20 ) );
BUF_X8 fanout_buf_21 ( .A(fanout_net_75 ), .Z(fanout_net_21 ) );
BUF_X8 fanout_buf_22 ( .A(fanout_net_75 ), .Z(fanout_net_22 ) );
BUF_X8 fanout_buf_23 ( .A(fanout_net_75 ), .Z(fanout_net_23 ) );
BUF_X8 fanout_buf_24 ( .A(fanout_net_75 ), .Z(fanout_net_24 ) );
BUF_X8 fanout_buf_25 ( .A(fanout_net_75 ), .Z(fanout_net_25 ) );
BUF_X8 fanout_buf_26 ( .A(fanout_net_75 ), .Z(fanout_net_26 ) );
BUF_X8 fanout_buf_27 ( .A(fanout_net_75 ), .Z(fanout_net_27 ) );
BUF_X8 fanout_buf_28 ( .A(fanout_net_75 ), .Z(fanout_net_28 ) );
BUF_X8 fanout_buf_29 ( .A(fanout_net_75 ), .Z(fanout_net_29 ) );
BUF_X8 fanout_buf_30 ( .A(fanout_net_75 ), .Z(fanout_net_30 ) );
BUF_X8 fanout_buf_31 ( .A(fanout_net_75 ), .Z(fanout_net_31 ) );
BUF_X8 fanout_buf_32 ( .A(fanout_net_76 ), .Z(fanout_net_32 ) );
BUF_X8 fanout_buf_33 ( .A(fanout_net_76 ), .Z(fanout_net_33 ) );
BUF_X8 fanout_buf_34 ( .A(fanout_net_76 ), .Z(fanout_net_34 ) );
BUF_X8 fanout_buf_35 ( .A(fanout_net_76 ), .Z(fanout_net_35 ) );
BUF_X8 fanout_buf_36 ( .A(fanout_net_76 ), .Z(fanout_net_36 ) );
BUF_X8 fanout_buf_37 ( .A(fanout_net_76 ), .Z(fanout_net_37 ) );
BUF_X8 fanout_buf_38 ( .A(fanout_net_76 ), .Z(fanout_net_38 ) );
BUF_X8 fanout_buf_39 ( .A(fanout_net_76 ), .Z(fanout_net_39 ) );
BUF_X8 fanout_buf_40 ( .A(fanout_net_76 ), .Z(fanout_net_40 ) );
BUF_X8 fanout_buf_41 ( .A(fanout_net_76 ), .Z(fanout_net_41 ) );
BUF_X8 fanout_buf_42 ( .A(fanout_net_76 ), .Z(fanout_net_42 ) );
BUF_X8 fanout_buf_43 ( .A(fanout_net_76 ), .Z(fanout_net_43 ) );
BUF_X8 fanout_buf_44 ( .A(fanout_net_76 ), .Z(fanout_net_44 ) );
BUF_X8 fanout_buf_45 ( .A(fanout_net_76 ), .Z(fanout_net_45 ) );
BUF_X8 fanout_buf_46 ( .A(fanout_net_76 ), .Z(fanout_net_46 ) );
BUF_X8 fanout_buf_47 ( .A(fanout_net_76 ), .Z(fanout_net_47 ) );
BUF_X8 fanout_buf_48 ( .A(fanout_net_76 ), .Z(fanout_net_48 ) );
BUF_X8 fanout_buf_49 ( .A(fanout_net_76 ), .Z(fanout_net_49 ) );
BUF_X8 fanout_buf_50 ( .A(fanout_net_76 ), .Z(fanout_net_50 ) );
BUF_X8 fanout_buf_51 ( .A(fanout_net_76 ), .Z(fanout_net_51 ) );
BUF_X8 fanout_buf_52 ( .A(fanout_net_76 ), .Z(fanout_net_52 ) );
BUF_X8 fanout_buf_53 ( .A(fanout_net_76 ), .Z(fanout_net_53 ) );
BUF_X8 fanout_buf_54 ( .A(fanout_net_76 ), .Z(fanout_net_54 ) );
BUF_X8 fanout_buf_55 ( .A(fanout_net_76 ), .Z(fanout_net_55 ) );
BUF_X8 fanout_buf_56 ( .A(fanout_net_76 ), .Z(fanout_net_56 ) );
BUF_X8 fanout_buf_57 ( .A(fanout_net_76 ), .Z(fanout_net_57 ) );
BUF_X8 fanout_buf_58 ( .A(fanout_net_76 ), .Z(fanout_net_58 ) );
BUF_X8 fanout_buf_59 ( .A(fanout_net_76 ), .Z(fanout_net_59 ) );
BUF_X8 fanout_buf_60 ( .A(fanout_net_76 ), .Z(fanout_net_60 ) );
BUF_X8 fanout_buf_61 ( .A(fanout_net_76 ), .Z(fanout_net_61 ) );
BUF_X8 fanout_buf_62 ( .A(reset ), .Z(fanout_net_62 ) );
BUF_X8 fanout_buf_63 ( .A(reset ), .Z(fanout_net_63 ) );
BUF_X8 fanout_buf_64 ( .A(reset ), .Z(fanout_net_64 ) );
BUF_X8 fanout_buf_65 ( .A(reset ), .Z(fanout_net_65 ) );
BUF_X8 fanout_buf_66 ( .A(reset ), .Z(fanout_net_66 ) );
BUF_X8 fanout_buf_67 ( .A(reset ), .Z(fanout_net_67 ) );
BUF_X8 fanout_buf_68 ( .A(reset ), .Z(fanout_net_68 ) );
BUF_X8 fanout_buf_69 ( .A(reset ), .Z(fanout_net_69 ) );
BUF_X8 fanout_buf_70 ( .A(reset ), .Z(fanout_net_70 ) );
BUF_X8 fanout_buf_71 ( .A(reset ), .Z(fanout_net_71 ) );
BUF_X8 fanout_buf_72 ( .A(reset ), .Z(fanout_net_72 ) );
BUF_X8 fanout_buf_73 ( .A(reset ), .Z(fanout_net_73 ) );
BUF_X8 fanout_buf_74 ( .A(reset ), .Z(fanout_net_74 ) );
BUF_X8 fanout_buf_75 ( .A(reset ), .Z(fanout_net_75 ) );
BUF_X8 fanout_buf_76 ( .A(reset ), .Z(fanout_net_76 ) );

endmodule
