//Generate the verilog at 2025-10-16T18:10:31 by iSTA.
module top (
clk,
gpr_we,
reset,
alu_result,
inst,
load_data,
pc,
wdata
);

input clk ;
output gpr_we ;
input reset ;
output [31:0] alu_result ;
output [31:0] inst ;
output [31:0] load_data ;
output [31:0] pc ;
output [31:0] wdata ;

wire _000_ ;
wire _001_ ;
wire _002_ ;
wire _003_ ;
wire _004_ ;
wire _005_ ;
wire _006_ ;
wire _007_ ;
wire _008_ ;
wire _009_ ;
wire _010_ ;
wire _011_ ;
wire _012_ ;
wire _013_ ;
wire _014_ ;
wire _015_ ;
wire _016_ ;
wire _017_ ;
wire _018_ ;
wire _019_ ;
wire _020_ ;
wire _021_ ;
wire _022_ ;
wire _023_ ;
wire _024_ ;
wire _025_ ;
wire _026_ ;
wire _027_ ;
wire _028_ ;
wire _029_ ;
wire _030_ ;
wire _031_ ;
wire _032_ ;
wire _033_ ;
wire _034_ ;
wire _035_ ;
wire _036_ ;
wire _037_ ;
wire _038_ ;
wire _039_ ;
wire _040_ ;
wire _041_ ;
wire _042_ ;
wire _043_ ;
wire _044_ ;
wire _045_ ;
wire _046_ ;
wire _047_ ;
wire _048_ ;
wire _049_ ;
wire _050_ ;
wire _051_ ;
wire _052_ ;
wire _053_ ;
wire _054_ ;
wire _055_ ;
wire _056_ ;
wire _057_ ;
wire _058_ ;
wire _059_ ;
wire _060_ ;
wire _061_ ;
wire _062_ ;
wire _063_ ;
wire _064_ ;
wire _065_ ;
wire _066_ ;
wire _067_ ;
wire _068_ ;
wire _069_ ;
wire _070_ ;
wire _071_ ;
wire _072_ ;
wire _073_ ;
wire _074_ ;
wire _075_ ;
wire _076_ ;
wire _077_ ;
wire _078_ ;
wire _079_ ;
wire _080_ ;
wire _081_ ;
wire _082_ ;
wire _083_ ;
wire _084_ ;
wire _085_ ;
wire _086_ ;
wire _087_ ;
wire _088_ ;
wire _089_ ;
wire _090_ ;
wire _091_ ;
wire _092_ ;
wire _093_ ;
wire _094_ ;
wire _095_ ;
wire _096_ ;
wire _097_ ;
wire _098_ ;
wire _099_ ;
wire _100_ ;
wire _101_ ;
wire _102_ ;
wire _103_ ;
wire _104_ ;
wire _105_ ;
wire _106_ ;
wire _107_ ;
wire _108_ ;
wire _109_ ;
wire _110_ ;
wire _111_ ;
wire _112_ ;
wire _113_ ;
wire _114_ ;
wire _115_ ;
wire _116_ ;
wire _117_ ;
wire _118_ ;
wire _119_ ;
wire _120_ ;
wire _121_ ;
wire _122_ ;
wire _123_ ;
wire _124_ ;
wire _125_ ;
wire _126_ ;
wire _127_ ;
wire _128_ ;
wire _129_ ;
wire _130_ ;
wire _131_ ;
wire _132_ ;
wire _133_ ;
wire _134_ ;
wire _135_ ;
wire clk ;
wire gpr_we ;
wire reset ;
wire \u_ifu.reset_sync ;
wire \alu_result[0] ;
wire \alu_result[1] ;
wire \alu_result[2] ;
wire \alu_result[3] ;
wire \alu_result[4] ;
wire \alu_result[5] ;
wire \alu_result[6] ;
wire \alu_result[7] ;
wire \alu_result[8] ;
wire \alu_result[9] ;
wire \alu_result[10] ;
wire \alu_result[11] ;
wire \alu_result[12] ;
wire \alu_result[13] ;
wire \alu_result[14] ;
wire \alu_result[15] ;
wire \alu_result[16] ;
wire \alu_result[17] ;
wire \alu_result[18] ;
wire \alu_result[19] ;
wire \alu_result[20] ;
wire \alu_result[21] ;
wire \alu_result[22] ;
wire \alu_result[23] ;
wire \alu_result[24] ;
wire \alu_result[25] ;
wire \alu_result[26] ;
wire \alu_result[27] ;
wire \alu_result[28] ;
wire \alu_result[29] ;
wire \alu_result[30] ;
wire \alu_result[31] ;
wire \inst[0] ;
wire \inst[1] ;
wire \inst[2] ;
wire \inst[3] ;
wire \inst[4] ;
wire \inst[5] ;
wire \inst[6] ;
wire \inst[7] ;
wire \inst[8] ;
wire \inst[9] ;
wire \inst[10] ;
wire \inst[11] ;
wire \inst[12] ;
wire \inst[13] ;
wire \inst[14] ;
wire \inst[15] ;
wire \inst[16] ;
wire \inst[17] ;
wire \inst[18] ;
wire \inst[19] ;
wire \inst[20] ;
wire \inst[21] ;
wire \inst[22] ;
wire \inst[23] ;
wire \inst[24] ;
wire \inst[25] ;
wire \inst[26] ;
wire \inst[27] ;
wire \inst[28] ;
wire \inst[29] ;
wire \inst[30] ;
wire \inst[31] ;
wire \load_data[0] ;
wire \load_data[1] ;
wire \load_data[2] ;
wire \load_data[3] ;
wire \load_data[4] ;
wire \load_data[5] ;
wire \load_data[6] ;
wire \load_data[7] ;
wire \load_data[8] ;
wire \load_data[9] ;
wire \load_data[10] ;
wire \load_data[11] ;
wire \load_data[12] ;
wire \load_data[13] ;
wire \load_data[14] ;
wire \load_data[15] ;
wire \load_data[16] ;
wire \load_data[17] ;
wire \load_data[18] ;
wire \load_data[19] ;
wire \load_data[20] ;
wire \load_data[21] ;
wire \load_data[22] ;
wire \load_data[23] ;
wire \load_data[24] ;
wire \load_data[25] ;
wire \load_data[26] ;
wire \load_data[27] ;
wire \load_data[28] ;
wire \load_data[29] ;
wire \load_data[30] ;
wire \load_data[31] ;
wire \pc[0] ;
wire \pc[1] ;
wire \pc[2] ;
wire \pc[3] ;
wire \pc[4] ;
wire \pc[5] ;
wire \pc[6] ;
wire \pc[7] ;
wire \pc[8] ;
wire \pc[9] ;
wire \pc[10] ;
wire \pc[11] ;
wire \pc[12] ;
wire \pc[13] ;
wire \pc[14] ;
wire \pc[15] ;
wire \pc[16] ;
wire \pc[17] ;
wire \pc[18] ;
wire \pc[19] ;
wire \pc[20] ;
wire \pc[21] ;
wire \pc[22] ;
wire \pc[23] ;
wire \pc[24] ;
wire \pc[25] ;
wire \pc[26] ;
wire \pc[27] ;
wire \pc[28] ;
wire \pc[29] ;
wire \pc[30] ;
wire \pc[31] ;
wire \snpc[0] ;
wire \snpc[1] ;
wire \snpc[2] ;
wire \wdata[0] ;
wire \wdata[1] ;
wire \wdata[2] ;
wire \wdata[3] ;
wire \wdata[4] ;
wire \wdata[5] ;
wire \wdata[6] ;
wire \wdata[7] ;
wire \wdata[8] ;
wire \wdata[9] ;
wire \wdata[10] ;
wire \wdata[11] ;
wire \wdata[12] ;
wire \wdata[13] ;
wire \wdata[14] ;
wire \wdata[15] ;
wire \wdata[16] ;
wire \wdata[17] ;
wire \wdata[18] ;
wire \wdata[19] ;
wire \wdata[20] ;
wire \wdata[21] ;
wire \wdata[22] ;
wire \wdata[23] ;
wire \wdata[24] ;
wire \wdata[25] ;
wire \wdata[26] ;
wire \wdata[27] ;
wire \wdata[28] ;
wire \wdata[29] ;
wire \wdata[30] ;
wire \wdata[31] ;

assign alu_result[0] = gpr_we ;
assign alu_result[0] = \alu_result[0] ;
assign alu_result[0] = \alu_result[1] ;
assign alu_result[0] = \alu_result[2] ;
assign alu_result[0] = \alu_result[3] ;
assign alu_result[0] = \alu_result[4] ;
assign alu_result[0] = \alu_result[5] ;
assign alu_result[0] = \alu_result[6] ;
assign alu_result[0] = \alu_result[7] ;
assign alu_result[0] = \alu_result[8] ;
assign alu_result[0] = \alu_result[9] ;
assign alu_result[0] = \alu_result[10] ;
assign alu_result[0] = \alu_result[11] ;
assign alu_result[0] = \alu_result[12] ;
assign alu_result[0] = \alu_result[13] ;
assign alu_result[0] = \alu_result[14] ;
assign alu_result[0] = \alu_result[15] ;
assign alu_result[0] = \alu_result[16] ;
assign alu_result[0] = \alu_result[17] ;
assign alu_result[0] = \alu_result[18] ;
assign alu_result[0] = \alu_result[19] ;
assign alu_result[0] = \alu_result[20] ;
assign alu_result[0] = \alu_result[21] ;
assign alu_result[0] = \alu_result[22] ;
assign alu_result[0] = \alu_result[23] ;
assign alu_result[0] = \alu_result[24] ;
assign alu_result[0] = \alu_result[25] ;
assign alu_result[0] = \alu_result[26] ;
assign alu_result[0] = \alu_result[27] ;
assign alu_result[0] = \alu_result[28] ;
assign alu_result[0] = \alu_result[29] ;
assign alu_result[0] = \alu_result[30] ;
assign alu_result[0] = \alu_result[31] ;
assign alu_result[0] = \load_data[0] ;
assign alu_result[0] = \load_data[1] ;
assign alu_result[0] = \load_data[2] ;
assign alu_result[0] = \load_data[3] ;
assign alu_result[0] = \load_data[4] ;
assign alu_result[0] = \load_data[5] ;
assign alu_result[0] = \load_data[6] ;
assign alu_result[0] = \load_data[7] ;
assign alu_result[0] = \load_data[8] ;
assign alu_result[0] = \load_data[9] ;
assign alu_result[0] = \load_data[10] ;
assign alu_result[0] = \load_data[11] ;
assign alu_result[0] = \load_data[12] ;
assign alu_result[0] = \load_data[13] ;
assign alu_result[0] = \load_data[14] ;
assign alu_result[0] = \load_data[15] ;
assign alu_result[0] = \load_data[16] ;
assign alu_result[0] = \load_data[17] ;
assign alu_result[0] = \load_data[18] ;
assign alu_result[0] = \load_data[19] ;
assign alu_result[0] = \load_data[20] ;
assign alu_result[0] = \load_data[21] ;
assign alu_result[0] = \load_data[22] ;
assign alu_result[0] = \load_data[23] ;
assign alu_result[0] = \load_data[24] ;
assign alu_result[0] = \load_data[25] ;
assign alu_result[0] = \load_data[26] ;
assign alu_result[0] = \load_data[27] ;
assign alu_result[0] = \load_data[28] ;
assign alu_result[0] = \load_data[29] ;
assign alu_result[0] = \load_data[30] ;
assign alu_result[0] = \load_data[31] ;
assign alu_result[0] = \pc[0] ;
assign alu_result[0] = \pc[1] ;
assign pc[2] = \pc[2] ;
assign pc[3] = \pc[3] ;
assign pc[4] = \pc[4] ;
assign pc[5] = \pc[5] ;
assign pc[6] = \pc[6] ;
assign pc[7] = \pc[7] ;
assign pc[8] = \pc[8] ;
assign pc[9] = \pc[9] ;
assign pc[10] = \pc[10] ;
assign pc[11] = \pc[11] ;
assign pc[12] = \pc[12] ;
assign pc[13] = \pc[13] ;
assign pc[14] = \pc[14] ;
assign pc[15] = \pc[15] ;
assign pc[16] = \pc[16] ;
assign pc[17] = \pc[17] ;
assign pc[18] = \pc[18] ;
assign pc[19] = \pc[19] ;
assign pc[20] = \pc[20] ;
assign pc[21] = \pc[21] ;
assign pc[22] = \pc[22] ;
assign pc[23] = \pc[23] ;
assign pc[24] = \pc[24] ;
assign pc[25] = \pc[25] ;
assign pc[26] = \pc[26] ;
assign pc[27] = \pc[27] ;
assign pc[28] = \pc[28] ;
assign pc[29] = \pc[29] ;
assign pc[30] = \pc[30] ;
assign pc[31] = \pc[31] ;
assign alu_result[0] = \wdata[0] ;
assign alu_result[0] = \wdata[1] ;
assign alu_result[0] = \wdata[2] ;
assign alu_result[0] = \wdata[3] ;
assign alu_result[0] = \wdata[4] ;
assign alu_result[0] = \wdata[5] ;
assign alu_result[0] = \wdata[6] ;
assign alu_result[0] = \wdata[7] ;
assign alu_result[0] = \wdata[8] ;
assign alu_result[0] = \wdata[9] ;
assign alu_result[0] = \wdata[10] ;
assign alu_result[0] = \wdata[11] ;
assign alu_result[0] = \wdata[12] ;
assign alu_result[0] = \wdata[13] ;
assign alu_result[0] = \wdata[14] ;
assign alu_result[0] = \wdata[15] ;
assign alu_result[0] = \wdata[16] ;
assign alu_result[0] = \wdata[17] ;
assign alu_result[0] = \wdata[18] ;
assign alu_result[0] = \wdata[19] ;
assign alu_result[0] = \wdata[20] ;
assign alu_result[0] = \wdata[21] ;
assign alu_result[0] = \wdata[22] ;
assign alu_result[0] = \wdata[23] ;
assign alu_result[0] = \wdata[24] ;
assign alu_result[0] = \wdata[25] ;
assign alu_result[0] = \wdata[26] ;
assign alu_result[0] = \wdata[27] ;
assign alu_result[0] = \wdata[28] ;
assign alu_result[0] = \wdata[29] ;
assign alu_result[0] = \wdata[30] ;
assign alu_result[0] = \wdata[31] ;

AND2_X4 _136_ ( .A1(\pc[3] ), .A2(\pc[2] ), .ZN(_074_ ) );
AND2_X4 _137_ ( .A1(_074_ ), .A2(\pc[4] ), .ZN(_075_ ) );
AND2_X4 _138_ ( .A1(_075_ ), .A2(\pc[5] ), .ZN(_076_ ) );
AND4_X1 _139_ ( .A1(\pc[8] ), .A2(\pc[7] ), .A3(\pc[6] ), .A4(\pc[9] ), .ZN(_077_ ) );
AND2_X4 _140_ ( .A1(_076_ ), .A2(_077_ ), .ZN(_078_ ) );
AND2_X4 _141_ ( .A1(\pc[10] ), .A2(\pc[11] ), .ZN(_079_ ) );
AND3_X1 _142_ ( .A1(_079_ ), .A2(\pc[13] ), .A3(\pc[12] ), .ZN(_080_ ) );
AND2_X1 _143_ ( .A1(\pc[15] ), .A2(\pc[14] ), .ZN(_081_ ) );
AND2_X1 _144_ ( .A1(\pc[16] ), .A2(\pc[17] ), .ZN(_082_ ) );
AND3_X1 _145_ ( .A1(_080_ ), .A2(_081_ ), .A3(_082_ ), .ZN(_083_ ) );
AND2_X4 _146_ ( .A1(_078_ ), .A2(_083_ ), .ZN(_084_ ) );
NAND3_X1 _147_ ( .A1(\pc[21] ), .A2(\pc[19] ), .A3(\pc[18] ), .ZN(_085_ ) );
INV_X1 _148_ ( .A(\pc[20] ), .ZN(_086_ ) );
NOR2_X1 _149_ ( .A1(_085_ ), .A2(_086_ ), .ZN(_087_ ) );
AND2_X1 _150_ ( .A1(\pc[23] ), .A2(\pc[22] ), .ZN(_088_ ) );
AND4_X1 _151_ ( .A1(\pc[24] ), .A2(_087_ ), .A3(\pc[25] ), .A4(_088_ ), .ZN(_089_ ) );
AND2_X4 _152_ ( .A1(_084_ ), .A2(_089_ ), .ZN(_090_ ) );
AND4_X1 _153_ ( .A1(\pc[28] ), .A2(\pc[27] ), .A3(\pc[26] ), .A4(\pc[29] ), .ZN(_091_ ) );
AND2_X4 _154_ ( .A1(_090_ ), .A2(_091_ ), .ZN(_092_ ) );
AND2_X1 _155_ ( .A1(_092_ ), .A2(\pc[30] ), .ZN(_093_ ) );
INV_X1 _156_ ( .A(\u_ifu.reset_sync ), .ZN(_094_ ) );
BUF_X4 _157_ ( .A(_094_ ), .Z(_095_ ) );
OAI21_X1 _158_ ( .A(_095_ ), .B1(_092_ ), .B2(\pc[30] ), .ZN(_096_ ) );
NOR2_X1 _159_ ( .A1(_093_ ), .A2(_096_ ), .ZN(_000_ ) );
AND2_X1 _160_ ( .A1(\pc[27] ), .A2(\pc[26] ), .ZN(_097_ ) );
AND2_X4 _161_ ( .A1(_090_ ), .A2(_097_ ), .ZN(_098_ ) );
AOI21_X1 _162_ ( .A(\pc[29] ), .B1(_098_ ), .B2(\pc[28] ), .ZN(_099_ ) );
NOR3_X1 _163_ ( .A1(_099_ ), .A2(\u_ifu.reset_sync ), .A3(_092_ ), .ZN(_001_ ) );
AND2_X1 _164_ ( .A1(_084_ ), .A2(\pc[18] ), .ZN(_100_ ) );
AND2_X1 _165_ ( .A1(_100_ ), .A2(\pc[19] ), .ZN(_101_ ) );
OAI21_X1 _166_ ( .A(_095_ ), .B1(_101_ ), .B2(\pc[20] ), .ZN(_102_ ) );
AND3_X1 _167_ ( .A1(_100_ ), .A2(\pc[20] ), .A3(\pc[19] ), .ZN(_103_ ) );
NOR2_X1 _168_ ( .A1(_102_ ), .A2(_103_ ), .ZN(_002_ ) );
AOI21_X1 _169_ ( .A(\pc[19] ), .B1(_084_ ), .B2(\pc[18] ), .ZN(_104_ ) );
NOR3_X1 _170_ ( .A1(_101_ ), .A2(_104_ ), .A3(\u_ifu.reset_sync ), .ZN(_003_ ) );
OAI21_X1 _171_ ( .A(_095_ ), .B1(_084_ ), .B2(\pc[18] ), .ZN(_105_ ) );
NOR2_X1 _172_ ( .A1(_100_ ), .A2(_105_ ), .ZN(_004_ ) );
AND2_X1 _173_ ( .A1(_078_ ), .A2(_080_ ), .ZN(_030_ ) );
AND2_X1 _174_ ( .A1(_030_ ), .A2(_081_ ), .ZN(_031_ ) );
AOI21_X1 _175_ ( .A(\pc[17] ), .B1(_031_ ), .B2(\pc[16] ), .ZN(_032_ ) );
AND4_X1 _176_ ( .A1(_078_ ), .A2(_080_ ), .A3(_081_ ), .A4(_082_ ), .ZN(_033_ ) );
NOR3_X1 _177_ ( .A1(_032_ ), .A2(\u_ifu.reset_sync ), .A3(_033_ ), .ZN(_005_ ) );
OAI21_X1 _178_ ( .A(_094_ ), .B1(_031_ ), .B2(\pc[16] ), .ZN(_034_ ) );
AND2_X4 _179_ ( .A1(_078_ ), .A2(_079_ ), .ZN(_035_ ) );
AND2_X1 _180_ ( .A1(_035_ ), .A2(\pc[12] ), .ZN(_036_ ) );
AND3_X1 _181_ ( .A1(_036_ ), .A2(\pc[13] ), .A3(_081_ ), .ZN(_037_ ) );
AOI21_X1 _182_ ( .A(_034_ ), .B1(_037_ ), .B2(\pc[16] ), .ZN(_006_ ) );
AOI21_X1 _183_ ( .A(\pc[15] ), .B1(_030_ ), .B2(\pc[14] ), .ZN(_038_ ) );
NOR3_X1 _184_ ( .A1(_031_ ), .A2(_038_ ), .A3(\u_ifu.reset_sync ), .ZN(_007_ ) );
AND3_X1 _185_ ( .A1(_036_ ), .A2(\pc[14] ), .A3(\pc[13] ), .ZN(_039_ ) );
OAI21_X1 _186_ ( .A(_095_ ), .B1(_030_ ), .B2(\pc[14] ), .ZN(_040_ ) );
NOR2_X1 _187_ ( .A1(_039_ ), .A2(_040_ ), .ZN(_008_ ) );
AND2_X1 _188_ ( .A1(_036_ ), .A2(\pc[13] ), .ZN(_041_ ) );
AOI21_X1 _189_ ( .A(\pc[13] ), .B1(_035_ ), .B2(\pc[12] ), .ZN(_042_ ) );
NOR3_X1 _190_ ( .A1(_041_ ), .A2(\u_ifu.reset_sync ), .A3(_042_ ), .ZN(_009_ ) );
OAI21_X1 _191_ ( .A(_095_ ), .B1(_035_ ), .B2(\pc[12] ), .ZN(_043_ ) );
NOR2_X1 _192_ ( .A1(_036_ ), .A2(_043_ ), .ZN(_010_ ) );
AOI21_X1 _193_ ( .A(\pc[11] ), .B1(_078_ ), .B2(\pc[10] ), .ZN(_044_ ) );
NOR3_X1 _194_ ( .A1(_035_ ), .A2(_044_ ), .A3(\u_ifu.reset_sync ), .ZN(_011_ ) );
AND2_X1 _195_ ( .A1(_098_ ), .A2(\pc[28] ), .ZN(_045_ ) );
OAI21_X1 _196_ ( .A(_095_ ), .B1(_098_ ), .B2(\pc[28] ), .ZN(_046_ ) );
NOR2_X1 _197_ ( .A1(_045_ ), .A2(_046_ ), .ZN(_012_ ) );
OAI21_X1 _198_ ( .A(_094_ ), .B1(_078_ ), .B2(\pc[10] ), .ZN(_047_ ) );
AOI21_X1 _199_ ( .A(_047_ ), .B1(\pc[10] ), .B2(_078_ ), .ZN(_013_ ) );
AND2_X1 _200_ ( .A1(_076_ ), .A2(\pc[6] ), .ZN(_048_ ) );
AND2_X1 _201_ ( .A1(_048_ ), .A2(\pc[7] ), .ZN(_049_ ) );
AOI21_X1 _202_ ( .A(\pc[9] ), .B1(_049_ ), .B2(\pc[8] ), .ZN(_050_ ) );
NOR3_X1 _203_ ( .A1(_050_ ), .A2(\u_ifu.reset_sync ), .A3(_078_ ), .ZN(_014_ ) );
OAI21_X1 _204_ ( .A(_094_ ), .B1(_049_ ), .B2(\pc[8] ), .ZN(_051_ ) );
AOI21_X1 _205_ ( .A(_051_ ), .B1(\pc[8] ), .B2(_049_ ), .ZN(_015_ ) );
AOI21_X1 _206_ ( .A(\pc[7] ), .B1(_076_ ), .B2(\pc[6] ), .ZN(_052_ ) );
NOR3_X1 _207_ ( .A1(_049_ ), .A2(\u_ifu.reset_sync ), .A3(_052_ ), .ZN(_016_ ) );
OAI21_X1 _208_ ( .A(_095_ ), .B1(_076_ ), .B2(\pc[6] ), .ZN(_053_ ) );
NOR2_X1 _209_ ( .A1(_048_ ), .A2(_053_ ), .ZN(_017_ ) );
AOI21_X1 _210_ ( .A(\pc[5] ), .B1(_074_ ), .B2(\pc[4] ), .ZN(_054_ ) );
NOR3_X1 _211_ ( .A1(_076_ ), .A2(\u_ifu.reset_sync ), .A3(_054_ ), .ZN(_018_ ) );
OAI21_X1 _212_ ( .A(_095_ ), .B1(_074_ ), .B2(\pc[4] ), .ZN(_055_ ) );
NOR2_X1 _213_ ( .A1(_075_ ), .A2(_055_ ), .ZN(_019_ ) );
NOR2_X1 _214_ ( .A1(\pc[3] ), .A2(\pc[2] ), .ZN(_056_ ) );
NOR3_X1 _215_ ( .A1(_074_ ), .A2(_056_ ), .A3(\u_ifu.reset_sync ), .ZN(_020_ ) );
AND2_X1 _216_ ( .A1(_095_ ), .A2(\snpc[2] ), .ZN(_021_ ) );
AOI21_X1 _217_ ( .A(\pc[27] ), .B1(_090_ ), .B2(\pc[26] ), .ZN(_057_ ) );
AND4_X1 _218_ ( .A1(\pc[27] ), .A2(_084_ ), .A3(\pc[26] ), .A4(_089_ ), .ZN(_058_ ) );
NOR3_X1 _219_ ( .A1(_057_ ), .A2(\u_ifu.reset_sync ), .A3(_058_ ), .ZN(_022_ ) );
AND2_X1 _220_ ( .A1(_090_ ), .A2(\pc[26] ), .ZN(_059_ ) );
OAI21_X1 _221_ ( .A(_094_ ), .B1(_090_ ), .B2(\pc[26] ), .ZN(_060_ ) );
NOR2_X1 _222_ ( .A1(_059_ ), .A2(_060_ ), .ZN(_023_ ) );
AND3_X1 _223_ ( .A1(_084_ ), .A2(_087_ ), .A3(_088_ ), .ZN(_061_ ) );
AOI21_X1 _224_ ( .A(\pc[25] ), .B1(_061_ ), .B2(\pc[24] ), .ZN(_062_ ) );
NOR3_X1 _225_ ( .A1(_062_ ), .A2(\u_ifu.reset_sync ), .A3(_090_ ), .ZN(_024_ ) );
OAI21_X1 _226_ ( .A(_094_ ), .B1(_061_ ), .B2(\pc[24] ), .ZN(_063_ ) );
AND2_X1 _227_ ( .A1(_084_ ), .A2(_087_ ), .ZN(_064_ ) );
AND2_X1 _228_ ( .A1(_064_ ), .A2(_088_ ), .ZN(_065_ ) );
AOI21_X1 _229_ ( .A(_063_ ), .B1(\pc[24] ), .B2(_065_ ), .ZN(_025_ ) );
AOI21_X1 _230_ ( .A(\pc[23] ), .B1(_064_ ), .B2(\pc[22] ), .ZN(_066_ ) );
NOR3_X1 _231_ ( .A1(_066_ ), .A2(\u_ifu.reset_sync ), .A3(_061_ ), .ZN(_026_ ) );
AND2_X1 _232_ ( .A1(_064_ ), .A2(\pc[22] ), .ZN(_067_ ) );
OAI21_X1 _233_ ( .A(_094_ ), .B1(_064_ ), .B2(\pc[22] ), .ZN(_068_ ) );
NOR2_X1 _234_ ( .A1(_067_ ), .A2(_068_ ), .ZN(_027_ ) );
NAND3_X1 _235_ ( .A1(_084_ ), .A2(\pc[19] ), .A3(\pc[18] ), .ZN(_069_ ) );
OR3_X2 _236_ ( .A1(_069_ ), .A2(\pc[21] ), .A3(_086_ ), .ZN(_070_ ) );
OAI21_X1 _237_ ( .A(\pc[21] ), .B1(_069_ ), .B2(_086_ ), .ZN(_071_ ) );
AOI21_X1 _238_ ( .A(\u_ifu.reset_sync ), .B1(_070_ ), .B2(_071_ ), .ZN(_028_ ) );
AOI21_X1 _239_ ( .A(\pc[31] ), .B1(_092_ ), .B2(\pc[30] ), .ZN(_072_ ) );
AND4_X1 _240_ ( .A1(\pc[30] ), .A2(_090_ ), .A3(\pc[31] ), .A4(_091_ ), .ZN(_073_ ) );
OAI21_X1 _241_ ( .A(_095_ ), .B1(_072_ ), .B2(_073_ ), .ZN(_029_ ) );
LOGIC0_X1 _242_ ( .Z(\alu_result[0] ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q ( .D(_000_ ), .CK(clk ), .Q(\pc[30] ), .QN(_134_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_1 ( .D(_001_ ), .CK(clk ), .Q(\pc[29] ), .QN(_133_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_10 ( .D(_002_ ), .CK(clk ), .Q(\pc[20] ), .QN(_132_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_11 ( .D(_003_ ), .CK(clk ), .Q(\pc[19] ), .QN(_131_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_12 ( .D(_004_ ), .CK(clk ), .Q(\pc[18] ), .QN(_130_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_13 ( .D(_005_ ), .CK(clk ), .Q(\pc[17] ), .QN(_129_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_14 ( .D(_006_ ), .CK(clk ), .Q(\pc[16] ), .QN(_128_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_15 ( .D(_007_ ), .CK(clk ), .Q(\pc[15] ), .QN(_127_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_16 ( .D(_008_ ), .CK(clk ), .Q(\pc[14] ), .QN(_126_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_17 ( .D(_009_ ), .CK(clk ), .Q(\pc[13] ), .QN(_125_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_18 ( .D(_010_ ), .CK(clk ), .Q(\pc[12] ), .QN(_124_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_19 ( .D(_011_ ), .CK(clk ), .Q(\pc[11] ), .QN(_123_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_2 ( .D(_012_ ), .CK(clk ), .Q(\pc[28] ), .QN(_122_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_20 ( .D(_013_ ), .CK(clk ), .Q(\pc[10] ), .QN(_121_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_21 ( .D(_014_ ), .CK(clk ), .Q(\pc[9] ), .QN(_120_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_22 ( .D(_015_ ), .CK(clk ), .Q(\pc[8] ), .QN(_119_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_23 ( .D(_016_ ), .CK(clk ), .Q(\pc[7] ), .QN(_118_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_24 ( .D(_017_ ), .CK(clk ), .Q(\pc[6] ), .QN(_117_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_25 ( .D(_018_ ), .CK(clk ), .Q(\pc[5] ), .QN(_116_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_26 ( .D(_019_ ), .CK(clk ), .Q(\pc[4] ), .QN(_115_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_27 ( .D(_020_ ), .CK(clk ), .Q(\pc[3] ), .QN(_114_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_28 ( .D(_021_ ), .CK(clk ), .Q(\pc[2] ), .QN(\snpc[2] ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_3 ( .D(_022_ ), .CK(clk ), .Q(\pc[27] ), .QN(_113_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_4 ( .D(_023_ ), .CK(clk ), .Q(\pc[26] ), .QN(_112_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_5 ( .D(_024_ ), .CK(clk ), .Q(\pc[25] ), .QN(_111_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_6 ( .D(_025_ ), .CK(clk ), .Q(\pc[24] ), .QN(_110_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_7 ( .D(_026_ ), .CK(clk ), .Q(\pc[23] ), .QN(_109_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_8 ( .D(_027_ ), .CK(clk ), .Q(\pc[22] ), .QN(_108_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP0__Q_9 ( .D(_028_ ), .CK(clk ), .Q(\pc[21] ), .QN(_107_ ) );
DFF_X1 \u_ifu.pc_$_SDFF_PP1__Q ( .D(_029_ ), .CK(clk ), .Q(\pc[31] ), .QN(_135_ ) );
DFF_X1 \u_ifu.reset_sync_$_DFF_P__Q ( .D(reset ), .CK(clk ), .Q(\u_ifu.reset_sync ), .QN(_106_ ) );

endmodule
