// import alu_pkg::*;

// 指令类型枚举
typedef enum logic [2:0] {
    TYPE_R,  // R型指令，寄存器间操作
    TYPE_I,  // I型指令，带有立即数和寄存器操作数
    TYPE_S,  // S型指令，存储指令
    TYPE_B,  // B型指令，分支指令
    TYPE_U,  // U型指令，带有高位立即数
    TYPE_J,  // J型指令，JAL跳转指令
    TYPE_N   // none，无操作数类型
} inst_t;

/* verilator lint_off DECLFILENAME */

module top (
    input clk,   // 时钟信号
    input reset  // 复位信号
    // input [31:0] inst,  // 输入指令
    // output logic [31:0] pc  // 程序计数器输出
);

    // IFU：负责 PC 和取指
    logic [31:0] ifu_raddr, snpc, jump_target;  // pc renamed to ifu_raddr, snpc, 跳转目标地址
    logic        jump_en;
    logic [31:0] ifu_rdata;  // 当前指令, inst renamed to ifu_rdata
    IFU u_ifu (
        .clk(clk),
        .reset(reset),
        .jump_target(jump_target),
        .jump_en(jump_en),
        .ifu_raddr(ifu_raddr),  // pc renamed
        .snpc(snpc),
        .ifu_rdata(ifu_rdata)  // inst renamed
    );

    // IDU：负责指令解码
    // 解码信号
    logic [6:0] opcode, funct7;
    logic [ 2:0] funct3;
    logic [31:0] imm;
    logic [4:0] rs1, rs2, rd;
    inst_t inst_type;
    IDU u_idu (
        .ifu_rdata(ifu_rdata),  // inst renamed
        .opcode(opcode),
        .funct3(funct3),
        .funct7(funct7),
        .rd(rd),
        .rs1(rs1),
        .rs2(rs2),
        .imm(imm),
        .inst_type(inst_type)
    );

    // GPR：通用寄存器组
    logic [31:0] gpr_rdata1, gpr_rdata2, gpr_wdata;  // 读寄存器组数据1、2，写寄存器数据, renamed
    logic gpr_we;
    GPR u_gpr (
        .clk(clk),
        .reset(reset),
        .gpr_we(gpr_we && (|rd)),  // we renamed
        .gpr_waddr(rd),  // waddr renamed
        .gpr_wdata(gpr_wdata),  // wdata renamed
        .gpr_raddr1(rs1),  // raddr1 renamed
        .gpr_raddr2(rs2),  // raddr2 renamed
        .gpr_rdata1(gpr_rdata1),  // rdata1 renamed
        .gpr_rdata2(gpr_rdata2)  // rdata2 renamed
    );

    // CSR：控制状态寄存器
    logic [3:0][31:0] csr_wdata, csr_rdata;  // CSR写数据，读数据
    logic [3:0] csr_we;
    CSR u_csr (
        .clk(clk),
        .reset(reset),
        .csr_we(csr_we),  // we renamed
        .csr_wdata(csr_wdata),  // din renamed
        .csr_rdata(csr_rdata)  // dout renamed
    );


    // EXU：负责根据控制信号来进行运算和跳转
    logic [31:0] alu_result;  // ALU计算结果
    logic [31:0] csr_read_data;  // CSR读取的数据
    EXU u_exu (
        .opcode       (opcode),
        .funct3       (funct3),
        .funct7       (funct7),
        .gpr_rdata1   (gpr_rdata1),  // src1 renamed
        .gpr_rdata2   (gpr_rdata2),  // src2 renamed
        .imm          (imm),
        .ifu_raddr    (ifu_raddr),  // pc renamed
        .snpc         (snpc),
        .inst_type    (inst_type),
        .csr_rdata    (csr_rdata),
        .alu_result   (alu_result),
        .jump_target  (jump_target),
        .jump_en      (jump_en),
        .csr_we       (csr_we),
        .csr_wdata    (csr_wdata),
        .csr_read_data(csr_read_data)
    );

    // LSU：负责加载和存储指令的内存访问
    logic [31:0] load_data;  // 加载数据
    LSU u_lsu (
        .clk       (clk),
        .inst_type (inst_type),
        .opcode    (opcode),
        .funct3    (funct3),
        .ifu_raddr (ifu_raddr),  // pc renamed
        .alu_result(alu_result),  // addr renamed
        .gpr_rdata2(gpr_rdata2),  // store_data renamed
        .load_data (load_data)
    );

    // WBU：负责写回GPR
    WBU u_wbu (
        .inst_type    (inst_type),
        .opcode       (opcode),
        .funct3       (funct3),
        .ifu_raddr    (ifu_raddr),  // pc renamed
        .snpc         (snpc),
        .alu_result   (alu_result),
        .load_data    (load_data),
        .csr_read_data(csr_read_data),
        .gpr_wdata    (gpr_wdata),  // wdata renamed
        .gpr_we       (gpr_we)
    );

endmodule

// IFU(Instruction Fetch Unit) 负责根据当前PC从存储器中取出一条指令
module IFU (
    input         clk,
    input         reset,
    input  [31:0] jump_target,
    input         jump_en,
    output logic [31:0] ifu_raddr,  // pc renamed
    output logic [31:0] snpc,
    output logic [31:0] ifu_rdata  // inst renamed
);
    localparam int RESET_PC = 32'h80000000;
    logic reset_sync;
    logic [31:0] dnpc;

    // DPI 接口：从内存读取指令并上报 instruction + next pc
    import "DPI-C" function int pmem_read_npc(input int raddr);
    import "DPI-C" function void update_inst_npc(
        input int inst,
        input int dnpc
    );

    // 同步复位信号（保留原逻辑）
    always_ff @(posedge clk) begin
        if (reset) reset_sync <= 1'b1;
        else reset_sync <= 1'b0;
    end

    // 读取当前 PC 指令并通知 DPI
    always_comb ifu_rdata = pmem_read_npc(ifu_raddr);  // inst and pc renamed
    always_comb update_inst_npc(ifu_rdata, dnpc);  // inst renamed

    // PC 寄存器更新
    always_ff @(posedge clk) begin
        if (reset_sync) ifu_raddr <= RESET_PC;  // pc renamed
        else ifu_raddr <= dnpc;  // pc renamed
    end

    // snpc / dnpc 选择逻辑
    assign snpc = ifu_raddr + 4;  // pc renamed
    assign dnpc = jump_en ? jump_target : snpc;
endmodule

// IDU(Instruction Decode Unit) 负责对当前指令进行译码, 准备执行阶段需要使用的数据和控制信号
module IDU (
    input [31:0] ifu_rdata,  // 输入指令, inst renamed
    output [6:0] opcode,  // 操作码
    output [2:0] funct3,  // 功能码
    output [6:0] funct7,  // 功能码扩展
    output [4:0] rd,  // 目的寄存器编号
    output [4:0] rs1,  // 源寄存器1编号
    output [4:0] rs2,  // 源寄存器2编号
    output logic [31:0] imm,  // 立即数
    output inst_t inst_type  // 指令类型输出
);
    assign opcode = ifu_rdata[6:0];  // inst renamed
    assign funct3 = ifu_rdata[14:12];  // inst renamed
    assign funct7 = ifu_rdata[31:25];  // inst renamed
    assign rd = ifu_rdata[11:7];  // inst renamed
    assign rs1 = ifu_rdata[19:15];  // inst renamed
    assign rs2 = ifu_rdata[24:20];  // inst renamed

    always_comb begin
        unique case (opcode)
            7'b0110011: inst_type = TYPE_R;  // 寄存器类型
            7'b0010011, 7'b0000011, 7'b1100111, 7'b1110011: inst_type = TYPE_I;  // 立即数类型
            7'b0100011: inst_type = TYPE_S;  // 存储类型
            7'b1100011: inst_type = TYPE_B;  // 分支类型
            7'b0110111, 7'b0010111: inst_type = TYPE_U;  // 上位立即数类型
            7'b1101111: inst_type = TYPE_J;  // 跳转类型
            default: inst_type = TYPE_N;  // 无操作数类型
        endcase
    end
    always_comb begin
        unique case (inst_type)
            TYPE_I: imm = {{20{ifu_rdata[31]}}, ifu_rdata[31:20]};  // 符号扩展I型立即数, inst renamed
            TYPE_S: imm = {{20{ifu_rdata[31]}}, ifu_rdata[31:25], ifu_rdata[11:7]};  // 符号扩展S型立即数, inst renamed
            TYPE_B:
            imm = {
                {19{ifu_rdata[31]}}, ifu_rdata[31], ifu_rdata[7], ifu_rdata[30:25], ifu_rdata[11:8], 1'b0
            };  // 符号扩展B型立即数, inst renamed
            TYPE_U: imm = {ifu_rdata[31:12], 12'b0};  // U型立即数（高20位）, inst renamed
            TYPE_J:
            imm = {
                {11{ifu_rdata[31]}}, ifu_rdata[31], ifu_rdata[19:12], ifu_rdata[20], ifu_rdata[30:21], 1'b0
            };  // 符号扩展J型立即数, inst renamed
            default: imm = 32'h0;
        endcase
    end
endmodule

// GPR(General Purpose Register) 负责通用寄存器的读写
module GPR (
    input clk,  // 时钟信号
    input reset,  // 复位信号
    input gpr_we,  // 写使能信号, we renamed
    input [4:0] gpr_waddr,  // 写寄存器地址, waddr renamed
    input [31:0] gpr_wdata,  // 写数据, wdata renamed
    input [4:0] gpr_raddr1,  // 读寄存器1地址, raddr1 renamed
    input [4:0] gpr_raddr2,  // 读寄存器2地址, raddr2 renamed
    output logic [31:0] gpr_rdata1,  // 读寄存器1数据, rdata1 renamed
    output logic [31:0] gpr_rdata2  // 读寄存器2数据, rdata2 renamed
);
    logic [31:0] regfile[32];  // 寄存器文件

    // import "DPI-C" function void output_gprs(input [31:0] gprs[]);
    // always_comb output_gprs(regfile);  // 输出寄存器状态到DPI-C

    always_ff @(posedge clk) begin
        if (reset) begin
            for (int i = 0; i < 32; i++) regfile[i] <= 32'h0;  // 复位时清零所有寄存器
        end else if (gpr_we) begin  // we renamed
            regfile[gpr_waddr] <= gpr_wdata;  // waddr and wdata renamed
        end
        // write_gpr_npc(waddr, wdata);  // 更新DPI-C接口寄存器
    end


    import "DPI-C" function void write_gpr_npc(
        input logic [ 4:0] idx,
        input logic [31:0] data
    );
    always_comb begin
        if (gpr_we) write_gpr_npc(gpr_waddr, gpr_wdata);  // we, waddr, wdata renamed
    end

    always_comb begin
        gpr_rdata1 = (gpr_raddr1 == 5'b0) ? 32'h0 : regfile[gpr_raddr1];  // rdata1 and raddr1 renamed
        gpr_rdata2 = (gpr_raddr2 == 5'b0) ? 32'h0 : regfile[gpr_raddr2];  // rdata2 and raddr2 renamed
    end
endmodule

// CSR(Control and Status Register) 负责控制和状态寄存器的读写
module CSR #(
    localparam int N = 4  // CSR寄存器数量
) (
    input clk,  // 时钟信号
    input reset,  // 复位信号
    input [N-1:0] csr_we,  // 写使能信号, we renamed
    input [N-1:0][31:0] csr_wdata,  // CSR寄存器地址, din renamed
    output logic [N-1:0][31:0] csr_rdata  // CSR寄存器数据输出, dout renamed
);
    always_ff @(posedge clk) begin
        if (reset) csr_rdata <= '0;  // 复位时清零所有CSR寄存器
        else begin
            for (int i = 0; i < N; i++) if (csr_we[i]) csr_rdata[i] <= csr_wdata[i];  // we, din, dout renamed
        end
    end

    import "DPI-C" function void write_csr_npc(
        input logic [ 1:0] idx,
        input logic [31:0] data
    );

    always_comb begin
        for (int i = 0; i < N; i++)
        if (csr_we[i]) write_csr_npc(i[1:0], csr_wdata[i]);  // we and din renamed
    end

endmodule

// typedef enum logic [11:0] {
//     CSR_MTVEC   = 12'h305,
//     CSR_MEPC    = 12'h341,
//     CSR_MSTATUS = 12'h300,
//     CSR_MCAUSE  = 12'h342
// } csr_addr_t;

// EXU(Execute Unit) 负责根据控制信号控制ALU, 对数据进行计算
module EXU (
    input         [ 6:0]       opcode,
    input         [ 2:0]       funct3,
    input         [ 6:0]       funct7,
    input         [31:0]       gpr_rdata1,  // src1 renamed
    input         [31:0]       gpr_rdata2,  // src2 renamed
    input         [31:0]       imm,
    input         [31:0]       ifu_raddr,  // pc renamed
    input         [31:0]       snpc,
    input  inst_t              inst_type,
    input   [ 3:0][31:0] csr_rdata,
    output logic  [31:0]       alu_result,
    output logic  [31:0]       jump_target,
    output logic               jump_en,
    output logic  [ 3:0]       csr_we,
    output logic  [ 3:0][31:0] csr_wdata,
    output logic  [31:0]       csr_read_data
);
    import "DPI-C" function void NPCINV(input int pc);
    import "DPI-C" function void NPCTRAP();

    logic [31:0] alu_a, alu_b;
    alu_op_t alu_op;

    alu #(
        .WIDTH(32)
    ) u_alu (
        .A(alu_a),
        .B(alu_b),
        .ALUop(alu_op),
        .Result(alu_result)
    );

    function automatic logic [1:0] csr_addr_to_idx(input logic [11:0] addr);
        unique case (addr)
            12'h305: return 2'd0;
            12'h341: return 2'd1;
            12'h300: return 2'd2;
            12'h342: return 2'd3;
            default: return 2'd0;
        endcase
    endfunction

    always_comb begin
        jump_target = 32'h0;
        jump_en     = 1'b0;
        unique case (inst_type)
            TYPE_I: begin
                alu_a = gpr_rdata1;  // src1 renamed
                alu_b = imm;
                if (opcode == 7'b1100111) begin  // JALR
                    jump_target = {alu_result[31:1], 1'b0};
                    jump_en     = 1'b1;
                end else if (opcode == 7'b1110011 && funct3 == 3'b000) begin  // SYSTEM
                    unique case (imm)
                        32'h0: begin
                            // ECALL
                            jump_target = csr_rdata[0];
                            jump_en     = 1'b1;
                        end
                        32'h302: begin
                            // MRET
                            jump_target = csr_rdata[1];
                            jump_en     = 1'b1;
                        end
                        default: ;
                    endcase
                end
            end
            TYPE_R: begin
                alu_a = gpr_rdata1;  // src1 renamed
                alu_b = gpr_rdata2;  // src2 renamed
            end
            TYPE_U: begin
                alu_a = (opcode == 7'b0110111) ? 32'h0 : ifu_raddr;  // pc renamed
                alu_b = imm;
            end
            TYPE_J: begin
                alu_a       = ifu_raddr;  // pc renamed
                alu_b       = imm;
                jump_target = alu_result;
                jump_en     = 1'b1;
            end
            TYPE_B: begin
                alu_a = ifu_raddr;  // pc renamed
                alu_b = imm;
                jump_target = alu_result;
                unique case (funct3)
                    3'b000:  jump_en = (gpr_rdata1 == gpr_rdata2);  // src1 and src2 renamed
                    3'b001:  jump_en = (gpr_rdata1 != gpr_rdata2);  // src1 and src2 renamed
                    3'b100:  jump_en = ($signed(gpr_rdata1) < $signed(gpr_rdata2));  // src1 and src2 renamed
                    3'b101:  jump_en = ($signed(gpr_rdata1) >= $signed(gpr_rdata2));  // src1 and src2 renamed
                    3'b110:  jump_en = (gpr_rdata1 < gpr_rdata2);  // src1 and src2 renamed
                    3'b111:  jump_en = (gpr_rdata1 >= gpr_rdata2);  // src1 and src2 renamed
                    default: jump_en = 1'b0;
                endcase
            end
            TYPE_S: begin
                alu_a = gpr_rdata1;  // src1 renamed
                alu_b = imm;
            end
            default: begin
                alu_a = gpr_rdata1;  // src1 renamed
                alu_b = gpr_rdata2;  // src2 renamed
            end
        endcase
    end

    always_comb begin
        alu_op = ALU_ADD;
        if (opcode == 7'b0010011 || opcode == 7'b0110011) begin
            unique case (funct3)
                3'b000: begin  // ADD/ADDI 或 SUB
                    if (inst_type == TYPE_R && funct7 == 7'b0100000) alu_op = ALU_SUB;
                end
                3'b001:  alu_op = ALU_SLL;  // SLLI/SLL
                3'b010:  alu_op = ALU_SLT;  // SLTI/SLT
                3'b011:  alu_op = ALU_SLTU;  // SLTIU/SLTU
                3'b100:  alu_op = ALU_XOR;  // XORI/XOR
                3'b101:  alu_op = (funct7[5] == 1'b1) ? ALU_SRA : ALU_SRL;  // SRAI/SRA 或 SRLI/SRL
                3'b110:  alu_op = ALU_OR;  // ORI/OR
                3'b111:  alu_op = ALU_AND;  // ANDI/AND
                default: alu_op = ALU_ADD;
            endcase
        end
    end


    wire [1:0] csr_idx = csr_addr_to_idx(imm[11:0]);  // CSR寄存器索引
    logic [31:0] mstatus_ecall, mstatus_mret;  // mstatus临时变量
    always_comb begin
        csr_we        = '0;
        csr_wdata     = '0;
        csr_read_data = 32'h0;

        mstatus_ecall = csr_rdata[2];
        mstatus_mret  = csr_rdata[2];
        if (inst_type == TYPE_I && opcode == 7'b1110011) begin
            // CSR指令执行
            unique case (funct3)
                3'b000: begin
                    if (imm == 32'h0) begin
                        // ECALL
                        csr_we               = 4'b1110;
                        csr_wdata[1]         = ifu_raddr;
                        csr_wdata[3]         = 32'd11;
                        mstatus_ecall[7]     = mstatus_ecall[3];
                        mstatus_ecall[3]     = 1'b0;
                        mstatus_ecall[12:11] = 2'b11;
                        csr_wdata[2]         = mstatus_ecall;
                    end else if (imm == 32'h302) begin
                        // MRET
                        csr_we[2]           = 1'b1;
                        mstatus_mret[3]     = mstatus_mret[7];
                        mstatus_mret[7]     = 1'b1;
                        mstatus_mret[12:11] = 2'b00;
                        csr_wdata[2]        = mstatus_mret;
                    end else if (imm == 32'h1) begin
                        // EBREAK
                        NPCTRAP();
                    end else begin
                        // 不支持的系统指令保持兼容旧行为
                        NPCINV(ifu_raddr);
                    end
                end
                3'b001: begin
                    // CSRRW
                    csr_we[csr_idx]    = 1'b1;
                    csr_wdata[csr_idx] = gpr_rdata1;  // src1 renamed
                end
                3'b010: begin
                    // CSRRR
                    csr_read_data = csr_rdata[csr_idx];
                end
                default: NPCINV(ifu_raddr);  // pc renamed
            endcase
        end
    end

endmodule

// LSU(Load Store Unit) 负责根据控制信号控制存储器, 从存储器中读出数据, 或将数据写入存储器
module LSU (
    input          clk,
    input  inst_t        inst_type,
    input   [ 6:0] opcode,
    input   [ 2:0] funct3,
    input   [31:0] ifu_raddr,  // pc renamed
    input   [31:0] alu_result,  // addr renamed
    input   [31:0] gpr_rdata2,  // store_data renamed
    output logic  [31:0] load_data
);
    import "DPI-C" function int pmem_read_npc(input int raddr);
    import "DPI-C" function void pmem_write_npc(
        input int  waddr,
        input int  wdata,
        input byte wmask
    );
    import "DPI-C" function void NPCINV(input int pc);

    int mem_rdata_raw;

    // 加载逻辑
    always_comb begin
        load_data     = 32'h0;
        mem_rdata_raw = 0;
        if (inst_type == TYPE_I && opcode == 7'b0000011) begin
            mem_rdata_raw = pmem_read_npc(alu_result);  // addr renamed
            unique case (funct3)
                3'b000: load_data = {{24{mem_rdata_raw[7]}}, mem_rdata_raw[7:0]};  // LB
                3'b010: load_data = mem_rdata_raw;  // LW
                3'b001: load_data = {{16{mem_rdata_raw[15]}}, mem_rdata_raw[15:0]};  // LH
                3'b101: load_data = {16'b0, mem_rdata_raw[15:0]};  // LHU
                3'b100: load_data = {24'b0, mem_rdata_raw[7:0]};  // LBU
                default: begin
                    load_data = 32'h0;
                    NPCINV(ifu_raddr);  // pc renamed
                end
            endcase
        end
    end

    // 存储逻辑
    always_comb begin
        if (inst_type == TYPE_S && opcode == 7'b0100011) begin
            unique case (funct3)
                3'b000:  pmem_write_npc(alu_result, gpr_rdata2, 8'h1);  // addr and store_data renamed
                3'b001:  pmem_write_npc(alu_result, gpr_rdata2, 8'h3);  // addr and store_data renamed
                3'b010:  pmem_write_npc(alu_result, gpr_rdata2, 8'hf);  // addr and store_data renamed
                default: ;  // 不支持的 store 类型保持兼容旧行为
            endcase
        end
    end
endmodule

// WBU(WriteBack Unit): 将数据写入寄存器
module WBU (
    input  inst_t        inst_type,
    input   [ 6:0] opcode,
    input   [ 2:0] funct3,
    input   [31:0] ifu_raddr,  // pc renamed
    input   [31:0] snpc,
    input   [31:0] alu_result,
    input   [31:0] load_data,
    input   [31:0] csr_read_data,
    output logic  [31:0] gpr_wdata,  // wdata renamed
    output logic         gpr_we
);
    import "DPI-C" function void NPCINV(input int pc);

    always_comb begin
        gpr_wdata  = 32'h0;  // wdata renamed
        gpr_we = 1'b0;

        unique case (inst_type)
            TYPE_I: begin
                if (opcode == 7'b1100111) begin
                    // JALR
                    gpr_wdata  = snpc;
                    gpr_we = 1'b1;
                end else if (opcode == 7'b0000011) begin
                    // Load指令: 写回内存数据
                    gpr_wdata  = load_data;
                    gpr_we = 1'b1;
                end else if (opcode == 7'b1110011) begin
                    // CSR指令: 写回CSR读值
                    if (funct3 == 3'b010) begin
                        gpr_wdata  = csr_read_data;
                        gpr_we = 1'b1;
                    end
                end else begin
                    // 其他I型指令(算术/逻辑): 写回ALU结果
                    unique case (funct3)
                        3'b000, 3'b001, 3'b010, 3'b011, 3'b100, 3'b101, 3'b110, 3'b111: begin
                            gpr_wdata  = alu_result;  // wdata renamed
                            gpr_we = 1'b1;
                        end
                        default: NPCINV(ifu_raddr);  // pc renamed
                    endcase
                end
            end
            TYPE_R: begin
                unique case (funct3)
                    3'b000, 3'b001, 3'b010, 3'b011, 3'b100, 3'b101, 3'b110, 3'b111: begin
                        gpr_wdata  = alu_result;  // wdata renamed
                        gpr_we = 1'b1;
                    end
                    default: NPCINV(ifu_raddr);  // pc renamed
                endcase
            end
            TYPE_U: begin
                gpr_wdata  = alu_result;  // wdata renamed
                gpr_we = 1'b1;
            end
            TYPE_J: begin
                // JAL
                gpr_wdata  = snpc;
                gpr_we = 1'b1;
            end
            default: ;  // TYPE_B / TYPE_S / TYPE_N 不写回寄存器
        endcase
    end
endmodule

