//Generate the verilog at 2025-05-07T19:17:28 by iSTA.
module top (
btn,
clk,
rst,
seg
);

input btn ;
input clk ;
input rst ;
output [13:0] seg ;

wire _000_ ;
wire _001_ ;
wire _002_ ;
wire _003_ ;
wire _004_ ;
wire _005_ ;
wire _006_ ;
wire _007_ ;
wire _008_ ;
wire _009_ ;
wire _010_ ;
wire _011_ ;
wire _012_ ;
wire _013_ ;
wire _014_ ;
wire _015_ ;
wire _016_ ;
wire _017_ ;
wire _018_ ;
wire _019_ ;
wire _020_ ;
wire _021_ ;
wire _022_ ;
wire _023_ ;
wire _024_ ;
wire _025_ ;
wire _026_ ;
wire _027_ ;
wire _028_ ;
wire _029_ ;
wire _030_ ;
wire _031_ ;
wire _032_ ;
wire _033_ ;
wire _034_ ;
wire _035_ ;
wire _036_ ;
wire _037_ ;
wire _038_ ;
wire _039_ ;
wire _040_ ;
wire _041_ ;
wire _042_ ;
wire _043_ ;
wire _044_ ;
wire _045_ ;
wire _046_ ;
wire _047_ ;
wire _048_ ;
wire _049_ ;
wire _050_ ;
wire _051_ ;
wire _052_ ;
wire _053_ ;
wire btn ;
wire btn_$_ANDNOT__A_Y ;
wire btn_reg ;
wire clk ;
wire rst ;
wire seg_$_MUX__Y_13_A_$_MUX__Y_A ;
wire seg_$_MUX__Y_13_B_$_ANDNOT__Y_B ;
wire seg_$_MUX__Y_6_A_$_MUX__Y_A ;
wire seg_$_MUX__Y_6_B_$_ANDNOT__Y_B ;
wire x_$_DFFE_PP0P__Q_D ;
wire \bcd7seg0.b[0] ;
wire \bcd7seg0.b[1] ;
wire \bcd7seg0.b[2] ;
wire \bcd7seg0.b[3] ;
wire \bcd7seg1.b[0] ;
wire \bcd7seg1.b[1] ;
wire \bcd7seg1.b[2] ;
wire \bcd7seg1.b[3] ;
wire \seg[0] ;
wire \seg[1] ;
wire \seg[2] ;
wire \seg[3] ;
wire \seg[4] ;
wire \seg[5] ;
wire \seg[6] ;
wire \seg[7] ;
wire \seg[8] ;
wire \seg[9] ;
wire \seg[10] ;
wire \seg[11] ;
wire \seg[12] ;
wire \seg[13] ;

assign seg[0] = \seg[0] ;
assign seg[1] = \seg[1] ;
assign seg[2] = \seg[2] ;
assign seg[3] = \seg[3] ;
assign seg[4] = \seg[4] ;
assign seg[5] = \seg[5] ;
assign seg[6] = \seg[6] ;
assign seg[7] = \seg[7] ;
assign seg[8] = \seg[8] ;
assign seg[9] = \seg[9] ;
assign seg[10] = \seg[10] ;
assign seg[11] = \seg[11] ;
assign seg[12] = \seg[12] ;
assign seg[13] = \seg[13] ;

INV_X1 _054_ ( .A(rst ), .ZN(_000_ ) );
INV_X1 _055_ ( .A(btn ), .ZN(_001_ ) );
NOR2_X1 _056_ ( .A1(_001_ ), .A2(btn_reg ), .ZN(btn_$_ANDNOT__A_Y ) );
AND2_X4 _057_ ( .A1(\bcd7seg0.b[1] ), .A2(\bcd7seg0.b[0] ), .ZN(_002_ ) );
INV_X32 _058_ ( .A(\bcd7seg0.b[0] ), .ZN(_003_ ) );
NOR2_X4 _059_ ( .A1(_003_ ), .A2(\bcd7seg0.b[1] ), .ZN(_004_ ) );
MUX2_X2 _060_ ( .A(_002_ ), .B(_004_ ), .S(\bcd7seg0.b[2] ), .Z(_005_ ) );
NOR2_X1 _061_ ( .A1(\bcd7seg0.b[1] ), .A2(\bcd7seg0.b[0] ), .ZN(_006_ ) );
INV_X2 _062_ ( .A(\bcd7seg0.b[2] ), .ZN(_007_ ) );
MUX2_X1 _063_ ( .A(_006_ ), .B(_004_ ), .S(_007_ ), .Z(_008_ ) );
INV_X1 _064_ ( .A(\bcd7seg0.b[3] ), .ZN(_009_ ) );
MUX2_X2 _065_ ( .A(_005_ ), .B(_008_ ), .S(_009_ ), .Z(\seg[6] ) );
OR3_X2 _066_ ( .A1(_002_ ), .A2(_006_ ), .A3(_007_ ), .ZN(_010_ ) );
NOR2_X1 _067_ ( .A1(\bcd7seg0.b[2] ), .A2(\bcd7seg0.b[0] ), .ZN(_011_ ) );
OAI21_X1 _068_ ( .A(\bcd7seg0.b[3] ), .B1(_003_ ), .B2(\bcd7seg0.b[1] ), .ZN(_012_ ) );
OAI22_X1 _069_ ( .A1(_010_ ), .A2(\bcd7seg0.b[3] ), .B1(_011_ ), .B2(_012_ ), .ZN(\seg[5] ) );
INV_X1 _070_ ( .A(\bcd7seg1.b[3] ), .ZN(_013_ ) );
INV_X1 _071_ ( .A(\bcd7seg1.b[0] ), .ZN(_014_ ) );
NOR3_X1 _072_ ( .A1(_014_ ), .A2(\bcd7seg1.b[2] ), .A3(\bcd7seg1.b[1] ), .ZN(_015_ ) );
INV_X1 _073_ ( .A(\bcd7seg1.b[2] ), .ZN(_016_ ) );
NOR3_X1 _074_ ( .A1(_016_ ), .A2(\bcd7seg1.b[0] ), .A3(\bcd7seg1.b[1] ), .ZN(_017_ ) );
OAI21_X1 _075_ ( .A(_013_ ), .B1(_015_ ), .B2(_017_ ), .ZN(_018_ ) );
AND2_X1 _076_ ( .A1(\bcd7seg1.b[0] ), .A2(\bcd7seg1.b[1] ), .ZN(_019_ ) );
NAND2_X1 _077_ ( .A1(_019_ ), .A2(\bcd7seg1.b[2] ), .ZN(_020_ ) );
AND2_X1 _078_ ( .A1(_014_ ), .A2(\bcd7seg1.b[1] ), .ZN(_021_ ) );
NAND2_X1 _079_ ( .A1(_021_ ), .A2(_016_ ), .ZN(_022_ ) );
OAI211_X1 _080_ ( .A(_018_ ), .B(_020_ ), .C1(_013_ ), .C2(_022_ ), .ZN(\seg[10] ) );
NOR2_X1 _081_ ( .A1(\bcd7seg1.b[2] ), .A2(\bcd7seg1.b[0] ), .ZN(_023_ ) );
OR3_X1 _082_ ( .A1(_021_ ), .A2(\bcd7seg1.b[3] ), .A3(_023_ ), .ZN(_024_ ) );
NOR2_X1 _083_ ( .A1(_014_ ), .A2(\bcd7seg1.b[1] ), .ZN(_025_ ) );
NAND3_X1 _084_ ( .A1(_025_ ), .A2(\bcd7seg1.b[3] ), .A3(seg_$_MUX__Y_13_B_$_ANDNOT__Y_B ), .ZN(_026_ ) );
NAND2_X1 _085_ ( .A1(_024_ ), .A2(_026_ ), .ZN(\seg[9] ) );
NAND3_X1 _086_ ( .A1(_025_ ), .A2(\bcd7seg1.b[3] ), .A3(\bcd7seg1.b[2] ), .ZN(_027_ ) );
AOI21_X1 _087_ ( .A(_016_ ), .B1(\bcd7seg1.b[0] ), .B2(\bcd7seg1.b[1] ), .ZN(_028_ ) );
OAI21_X1 _088_ ( .A(_013_ ), .B1(\bcd7seg1.b[0] ), .B2(\bcd7seg1.b[1] ), .ZN(_029_ ) );
OAI21_X1 _089_ ( .A(_027_ ), .B1(_028_ ), .B2(_029_ ), .ZN(\seg[8] ) );
OR4_X4 _090_ ( .A1(_013_ ), .A2(\bcd7seg1.b[0] ), .A3(\bcd7seg1.b[1] ), .A4(seg_$_MUX__Y_13_B_$_ANDNOT__Y_B ), .ZN(_030_ ) );
OAI21_X1 _091_ ( .A(_013_ ), .B1(\bcd7seg1.b[2] ), .B2(seg_$_MUX__Y_13_A_$_MUX__Y_A ), .ZN(_031_ ) );
OAI21_X1 _092_ ( .A(_030_ ), .B1(_028_ ), .B2(_031_ ), .ZN(\seg[7] ) );
NAND3_X1 _093_ ( .A1(_011_ ), .A2(_009_ ), .A3(\bcd7seg0.b[1] ), .ZN(_032_ ) );
AOI22_X1 _094_ ( .A1(_032_ ), .A2(_012_ ), .B1(\bcd7seg0.b[3] ), .B2(_007_ ), .ZN(\seg[4] ) );
OAI211_X1 _095_ ( .A(_010_ ), .B(_009_ ), .C1(\bcd7seg0.b[2] ), .C2(_004_ ), .ZN(_033_ ) );
AOI22_X1 _096_ ( .A1(\bcd7seg0.b[2] ), .A2(_002_ ), .B1(_011_ ), .B2(\bcd7seg0.b[1] ), .ZN(_034_ ) );
OAI21_X1 _097_ ( .A(_033_ ), .B1(_009_ ), .B2(_034_ ), .ZN(\seg[3] ) );
OAI21_X1 _098_ ( .A(_003_ ), .B1(_007_ ), .B2(\bcd7seg0.b[1] ), .ZN(_035_ ) );
AND2_X1 _099_ ( .A1(_004_ ), .A2(seg_$_MUX__Y_6_B_$_ANDNOT__Y_B ), .ZN(_036_ ) );
MUX2_X1 _100_ ( .A(_035_ ), .B(_036_ ), .S(\bcd7seg0.b[3] ), .Z(\seg[2] ) );
AND2_X1 _101_ ( .A1(_002_ ), .A2(\bcd7seg0.b[2] ), .ZN(_037_ ) );
NOR2_X1 _102_ ( .A1(_006_ ), .A2(\bcd7seg0.b[2] ), .ZN(_038_ ) );
OAI21_X1 _103_ ( .A(_009_ ), .B1(_037_ ), .B2(_038_ ), .ZN(_039_ ) );
NAND3_X1 _104_ ( .A1(_004_ ), .A2(\bcd7seg0.b[3] ), .A3(\bcd7seg0.b[2] ), .ZN(_040_ ) );
NAND2_X1 _105_ ( .A1(_039_ ), .A2(_040_ ), .ZN(\seg[1] ) );
OR4_X4 _106_ ( .A1(_009_ ), .A2(\bcd7seg0.b[1] ), .A3(\bcd7seg0.b[0] ), .A4(seg_$_MUX__Y_6_B_$_ANDNOT__Y_B ), .ZN(_041_ ) );
AOI21_X1 _107_ ( .A(_037_ ), .B1(_007_ ), .B2(seg_$_MUX__Y_6_A_$_MUX__Y_A ), .ZN(_042_ ) );
OAI21_X1 _108_ ( .A(_041_ ), .B1(_042_ ), .B2(\bcd7seg0.b[3] ), .ZN(\seg[0] ) );
NAND3_X1 _109_ ( .A1(_019_ ), .A2(\bcd7seg1.b[3] ), .A3(_016_ ), .ZN(_043_ ) );
NAND3_X1 _110_ ( .A1(_018_ ), .A2(_027_ ), .A3(_043_ ), .ZN(\seg[13] ) );
OAI211_X1 _111_ ( .A(_028_ ), .B(_013_ ), .C1(\bcd7seg1.b[0] ), .C2(\bcd7seg1.b[1] ), .ZN(_044_ ) );
OAI21_X1 _112_ ( .A(\bcd7seg1.b[3] ), .B1(_014_ ), .B2(\bcd7seg1.b[1] ), .ZN(_045_ ) );
OAI21_X1 _113_ ( .A(_044_ ), .B1(_023_ ), .B2(_045_ ), .ZN(\seg[12] ) );
AOI22_X1 _114_ ( .A1(_022_ ), .A2(_045_ ), .B1(\bcd7seg1.b[3] ), .B2(_016_ ), .ZN(\seg[11] ) );
XNOR2_X1 _115_ ( .A(\bcd7seg0.b[3] ), .B(\bcd7seg1.b[0] ), .ZN(_046_ ) );
XNOR2_X1 _116_ ( .A(\bcd7seg0.b[0] ), .B(seg_$_MUX__Y_6_B_$_ANDNOT__Y_B ), .ZN(_047_ ) );
XNOR2_X1 _117_ ( .A(_046_ ), .B(_047_ ), .ZN(x_$_DFFE_PP0P__Q_D ) );
CLKGATE_X1 _118_ ( .CK(clk ), .E(btn_$_ANDNOT__A_Y ), .GCK(_048_ ) );
DFFR_X1 btn_reg_$_DFF_PP0__Q ( .D(btn ), .RN(_000_ ), .CK(clk ), .Q(btn_reg ), .QN(_052_ ) );
DFFR_X1 x_$_DFFE_PP0P__Q ( .D(x_$_DFFE_PP0P__Q_D ), .RN(_000_ ), .CK(_048_ ), .Q(\bcd7seg1.b[3] ), .QN(_053_ ) );
DFFR_X1 x_$_DFFE_PP0P__Q_1 ( .D(\bcd7seg1.b[3] ), .RN(_000_ ), .CK(_048_ ), .Q(\bcd7seg1.b[2] ), .QN(seg_$_MUX__Y_13_B_$_ANDNOT__Y_B ) );
DFFR_X1 x_$_DFFE_PP0P__Q_2 ( .D(\bcd7seg1.b[2] ), .RN(_000_ ), .CK(_048_ ), .Q(\bcd7seg1.b[1] ), .QN(seg_$_MUX__Y_13_A_$_MUX__Y_A ) );
DFFR_X1 x_$_DFFE_PP0P__Q_3 ( .D(\bcd7seg1.b[1] ), .RN(_000_ ), .CK(_048_ ), .Q(\bcd7seg1.b[0] ), .QN(_051_ ) );
DFFR_X1 x_$_DFFE_PP0P__Q_4 ( .D(\bcd7seg1.b[0] ), .RN(_000_ ), .CK(_048_ ), .Q(\bcd7seg0.b[3] ), .QN(_050_ ) );
DFFR_X1 x_$_DFFE_PP0P__Q_5 ( .D(\bcd7seg0.b[3] ), .RN(_000_ ), .CK(_048_ ), .Q(\bcd7seg0.b[2] ), .QN(seg_$_MUX__Y_6_B_$_ANDNOT__Y_B ) );
DFFR_X1 x_$_DFFE_PP0P__Q_6 ( .D(\bcd7seg0.b[2] ), .RN(_000_ ), .CK(_048_ ), .Q(\bcd7seg0.b[1] ), .QN(seg_$_MUX__Y_6_A_$_MUX__Y_A ) );
DFFS_X1 x_$_DFFE_PP1P__Q ( .D(\bcd7seg0.b[1] ), .SN(_000_ ), .CK(_048_ ), .Q(\bcd7seg0.b[0] ), .QN(_049_ ) );

endmodule
